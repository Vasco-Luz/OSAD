magic
tech sky130A
magscale 1 2
timestamp 1743851084
<< pwell >>
rect -26 -26 12646 226
<< nmos >>
rect 60 0 860 200
rect 960 0 1760 200
rect 1860 0 2660 200
rect 2760 0 3560 200
rect 3660 0 4460 200
rect 4560 0 5360 200
rect 5460 0 6260 200
rect 6360 0 7160 200
rect 7260 0 8060 200
rect 8160 0 8960 200
rect 9060 0 9860 200
rect 9960 0 10760 200
rect 10860 0 11660 200
rect 11760 0 12560 200
<< ndiff >>
rect 0 153 60 200
rect 0 119 13 153
rect 47 119 60 153
rect 0 81 60 119
rect 0 47 13 81
rect 47 47 60 81
rect 0 0 60 47
rect 860 153 960 200
rect 860 119 893 153
rect 927 119 960 153
rect 860 81 960 119
rect 860 47 893 81
rect 927 47 960 81
rect 860 0 960 47
rect 1760 153 1860 200
rect 1760 119 1793 153
rect 1827 119 1860 153
rect 1760 81 1860 119
rect 1760 47 1793 81
rect 1827 47 1860 81
rect 1760 0 1860 47
rect 2660 153 2760 200
rect 2660 119 2693 153
rect 2727 119 2760 153
rect 2660 81 2760 119
rect 2660 47 2693 81
rect 2727 47 2760 81
rect 2660 0 2760 47
rect 3560 153 3660 200
rect 3560 119 3593 153
rect 3627 119 3660 153
rect 3560 81 3660 119
rect 3560 47 3593 81
rect 3627 47 3660 81
rect 3560 0 3660 47
rect 4460 153 4560 200
rect 4460 119 4493 153
rect 4527 119 4560 153
rect 4460 81 4560 119
rect 4460 47 4493 81
rect 4527 47 4560 81
rect 4460 0 4560 47
rect 5360 153 5460 200
rect 5360 119 5393 153
rect 5427 119 5460 153
rect 5360 81 5460 119
rect 5360 47 5393 81
rect 5427 47 5460 81
rect 5360 0 5460 47
rect 6260 153 6360 200
rect 6260 119 6293 153
rect 6327 119 6360 153
rect 6260 81 6360 119
rect 6260 47 6293 81
rect 6327 47 6360 81
rect 6260 0 6360 47
rect 7160 153 7260 200
rect 7160 119 7193 153
rect 7227 119 7260 153
rect 7160 81 7260 119
rect 7160 47 7193 81
rect 7227 47 7260 81
rect 7160 0 7260 47
rect 8060 153 8160 200
rect 8060 119 8093 153
rect 8127 119 8160 153
rect 8060 81 8160 119
rect 8060 47 8093 81
rect 8127 47 8160 81
rect 8060 0 8160 47
rect 8960 153 9060 200
rect 8960 119 8993 153
rect 9027 119 9060 153
rect 8960 81 9060 119
rect 8960 47 8993 81
rect 9027 47 9060 81
rect 8960 0 9060 47
rect 9860 153 9960 200
rect 9860 119 9893 153
rect 9927 119 9960 153
rect 9860 81 9960 119
rect 9860 47 9893 81
rect 9927 47 9960 81
rect 9860 0 9960 47
rect 10760 153 10860 200
rect 10760 119 10793 153
rect 10827 119 10860 153
rect 10760 81 10860 119
rect 10760 47 10793 81
rect 10827 47 10860 81
rect 10760 0 10860 47
rect 11660 153 11760 200
rect 11660 119 11693 153
rect 11727 119 11760 153
rect 11660 81 11760 119
rect 11660 47 11693 81
rect 11727 47 11760 81
rect 11660 0 11760 47
rect 12560 153 12620 200
rect 12560 119 12573 153
rect 12607 119 12620 153
rect 12560 81 12620 119
rect 12560 47 12573 81
rect 12607 47 12620 81
rect 12560 0 12620 47
<< ndiffc >>
rect 13 119 47 153
rect 13 47 47 81
rect 893 119 927 153
rect 893 47 927 81
rect 1793 119 1827 153
rect 1793 47 1827 81
rect 2693 119 2727 153
rect 2693 47 2727 81
rect 3593 119 3627 153
rect 3593 47 3627 81
rect 4493 119 4527 153
rect 4493 47 4527 81
rect 5393 119 5427 153
rect 5393 47 5427 81
rect 6293 119 6327 153
rect 6293 47 6327 81
rect 7193 119 7227 153
rect 7193 47 7227 81
rect 8093 119 8127 153
rect 8093 47 8127 81
rect 8993 119 9027 153
rect 8993 47 9027 81
rect 9893 119 9927 153
rect 9893 47 9927 81
rect 10793 119 10827 153
rect 10793 47 10827 81
rect 11693 119 11727 153
rect 11693 47 11727 81
rect 12573 119 12607 153
rect 12573 47 12607 81
<< poly >>
rect 60 290 860 306
rect 60 256 83 290
rect 117 256 155 290
rect 189 256 227 290
rect 261 256 299 290
rect 333 256 371 290
rect 405 256 443 290
rect 477 256 515 290
rect 549 256 587 290
rect 621 256 659 290
rect 693 256 731 290
rect 765 256 803 290
rect 837 256 860 290
rect 60 200 860 256
rect 960 290 1760 306
rect 960 256 983 290
rect 1017 256 1055 290
rect 1089 256 1127 290
rect 1161 256 1199 290
rect 1233 256 1271 290
rect 1305 256 1343 290
rect 1377 256 1415 290
rect 1449 256 1487 290
rect 1521 256 1559 290
rect 1593 256 1631 290
rect 1665 256 1703 290
rect 1737 256 1760 290
rect 960 200 1760 256
rect 1860 290 2660 306
rect 1860 256 1883 290
rect 1917 256 1955 290
rect 1989 256 2027 290
rect 2061 256 2099 290
rect 2133 256 2171 290
rect 2205 256 2243 290
rect 2277 256 2315 290
rect 2349 256 2387 290
rect 2421 256 2459 290
rect 2493 256 2531 290
rect 2565 256 2603 290
rect 2637 256 2660 290
rect 1860 200 2660 256
rect 2760 290 3560 306
rect 2760 256 2783 290
rect 2817 256 2855 290
rect 2889 256 2927 290
rect 2961 256 2999 290
rect 3033 256 3071 290
rect 3105 256 3143 290
rect 3177 256 3215 290
rect 3249 256 3287 290
rect 3321 256 3359 290
rect 3393 256 3431 290
rect 3465 256 3503 290
rect 3537 256 3560 290
rect 2760 200 3560 256
rect 3660 290 4460 306
rect 3660 256 3683 290
rect 3717 256 3755 290
rect 3789 256 3827 290
rect 3861 256 3899 290
rect 3933 256 3971 290
rect 4005 256 4043 290
rect 4077 256 4115 290
rect 4149 256 4187 290
rect 4221 256 4259 290
rect 4293 256 4331 290
rect 4365 256 4403 290
rect 4437 256 4460 290
rect 3660 200 4460 256
rect 4560 290 5360 306
rect 4560 256 4583 290
rect 4617 256 4655 290
rect 4689 256 4727 290
rect 4761 256 4799 290
rect 4833 256 4871 290
rect 4905 256 4943 290
rect 4977 256 5015 290
rect 5049 256 5087 290
rect 5121 256 5159 290
rect 5193 256 5231 290
rect 5265 256 5303 290
rect 5337 256 5360 290
rect 4560 200 5360 256
rect 5460 290 6260 306
rect 5460 256 5483 290
rect 5517 256 5555 290
rect 5589 256 5627 290
rect 5661 256 5699 290
rect 5733 256 5771 290
rect 5805 256 5843 290
rect 5877 256 5915 290
rect 5949 256 5987 290
rect 6021 256 6059 290
rect 6093 256 6131 290
rect 6165 256 6203 290
rect 6237 256 6260 290
rect 5460 200 6260 256
rect 6360 290 7160 306
rect 6360 256 6383 290
rect 6417 256 6455 290
rect 6489 256 6527 290
rect 6561 256 6599 290
rect 6633 256 6671 290
rect 6705 256 6743 290
rect 6777 256 6815 290
rect 6849 256 6887 290
rect 6921 256 6959 290
rect 6993 256 7031 290
rect 7065 256 7103 290
rect 7137 256 7160 290
rect 6360 200 7160 256
rect 7260 290 8060 306
rect 7260 256 7283 290
rect 7317 256 7355 290
rect 7389 256 7427 290
rect 7461 256 7499 290
rect 7533 256 7571 290
rect 7605 256 7643 290
rect 7677 256 7715 290
rect 7749 256 7787 290
rect 7821 256 7859 290
rect 7893 256 7931 290
rect 7965 256 8003 290
rect 8037 256 8060 290
rect 7260 200 8060 256
rect 8160 290 8960 306
rect 8160 256 8183 290
rect 8217 256 8255 290
rect 8289 256 8327 290
rect 8361 256 8399 290
rect 8433 256 8471 290
rect 8505 256 8543 290
rect 8577 256 8615 290
rect 8649 256 8687 290
rect 8721 256 8759 290
rect 8793 256 8831 290
rect 8865 256 8903 290
rect 8937 256 8960 290
rect 8160 200 8960 256
rect 9060 290 9860 306
rect 9060 256 9083 290
rect 9117 256 9155 290
rect 9189 256 9227 290
rect 9261 256 9299 290
rect 9333 256 9371 290
rect 9405 256 9443 290
rect 9477 256 9515 290
rect 9549 256 9587 290
rect 9621 256 9659 290
rect 9693 256 9731 290
rect 9765 256 9803 290
rect 9837 256 9860 290
rect 9060 200 9860 256
rect 9960 290 10760 306
rect 9960 256 9983 290
rect 10017 256 10055 290
rect 10089 256 10127 290
rect 10161 256 10199 290
rect 10233 256 10271 290
rect 10305 256 10343 290
rect 10377 256 10415 290
rect 10449 256 10487 290
rect 10521 256 10559 290
rect 10593 256 10631 290
rect 10665 256 10703 290
rect 10737 256 10760 290
rect 9960 200 10760 256
rect 10860 290 11660 306
rect 10860 256 10883 290
rect 10917 256 10955 290
rect 10989 256 11027 290
rect 11061 256 11099 290
rect 11133 256 11171 290
rect 11205 256 11243 290
rect 11277 256 11315 290
rect 11349 256 11387 290
rect 11421 256 11459 290
rect 11493 256 11531 290
rect 11565 256 11603 290
rect 11637 256 11660 290
rect 10860 200 11660 256
rect 11760 290 12560 306
rect 11760 256 11783 290
rect 11817 256 11855 290
rect 11889 256 11927 290
rect 11961 256 11999 290
rect 12033 256 12071 290
rect 12105 256 12143 290
rect 12177 256 12215 290
rect 12249 256 12287 290
rect 12321 256 12359 290
rect 12393 256 12431 290
rect 12465 256 12503 290
rect 12537 256 12560 290
rect 11760 200 12560 256
rect 60 -40 860 0
rect 960 -40 1760 0
rect 1860 -40 2660 0
rect 2760 -40 3560 0
rect 3660 -40 4460 0
rect 4560 -40 5360 0
rect 5460 -40 6260 0
rect 6360 -40 7160 0
rect 7260 -40 8060 0
rect 8160 -40 8960 0
rect 9060 -40 9860 0
rect 9960 -40 10760 0
rect 10860 -40 11660 0
rect 11760 -40 12560 0
<< polycont >>
rect 83 256 117 290
rect 155 256 189 290
rect 227 256 261 290
rect 299 256 333 290
rect 371 256 405 290
rect 443 256 477 290
rect 515 256 549 290
rect 587 256 621 290
rect 659 256 693 290
rect 731 256 765 290
rect 803 256 837 290
rect 983 256 1017 290
rect 1055 256 1089 290
rect 1127 256 1161 290
rect 1199 256 1233 290
rect 1271 256 1305 290
rect 1343 256 1377 290
rect 1415 256 1449 290
rect 1487 256 1521 290
rect 1559 256 1593 290
rect 1631 256 1665 290
rect 1703 256 1737 290
rect 1883 256 1917 290
rect 1955 256 1989 290
rect 2027 256 2061 290
rect 2099 256 2133 290
rect 2171 256 2205 290
rect 2243 256 2277 290
rect 2315 256 2349 290
rect 2387 256 2421 290
rect 2459 256 2493 290
rect 2531 256 2565 290
rect 2603 256 2637 290
rect 2783 256 2817 290
rect 2855 256 2889 290
rect 2927 256 2961 290
rect 2999 256 3033 290
rect 3071 256 3105 290
rect 3143 256 3177 290
rect 3215 256 3249 290
rect 3287 256 3321 290
rect 3359 256 3393 290
rect 3431 256 3465 290
rect 3503 256 3537 290
rect 3683 256 3717 290
rect 3755 256 3789 290
rect 3827 256 3861 290
rect 3899 256 3933 290
rect 3971 256 4005 290
rect 4043 256 4077 290
rect 4115 256 4149 290
rect 4187 256 4221 290
rect 4259 256 4293 290
rect 4331 256 4365 290
rect 4403 256 4437 290
rect 4583 256 4617 290
rect 4655 256 4689 290
rect 4727 256 4761 290
rect 4799 256 4833 290
rect 4871 256 4905 290
rect 4943 256 4977 290
rect 5015 256 5049 290
rect 5087 256 5121 290
rect 5159 256 5193 290
rect 5231 256 5265 290
rect 5303 256 5337 290
rect 5483 256 5517 290
rect 5555 256 5589 290
rect 5627 256 5661 290
rect 5699 256 5733 290
rect 5771 256 5805 290
rect 5843 256 5877 290
rect 5915 256 5949 290
rect 5987 256 6021 290
rect 6059 256 6093 290
rect 6131 256 6165 290
rect 6203 256 6237 290
rect 6383 256 6417 290
rect 6455 256 6489 290
rect 6527 256 6561 290
rect 6599 256 6633 290
rect 6671 256 6705 290
rect 6743 256 6777 290
rect 6815 256 6849 290
rect 6887 256 6921 290
rect 6959 256 6993 290
rect 7031 256 7065 290
rect 7103 256 7137 290
rect 7283 256 7317 290
rect 7355 256 7389 290
rect 7427 256 7461 290
rect 7499 256 7533 290
rect 7571 256 7605 290
rect 7643 256 7677 290
rect 7715 256 7749 290
rect 7787 256 7821 290
rect 7859 256 7893 290
rect 7931 256 7965 290
rect 8003 256 8037 290
rect 8183 256 8217 290
rect 8255 256 8289 290
rect 8327 256 8361 290
rect 8399 256 8433 290
rect 8471 256 8505 290
rect 8543 256 8577 290
rect 8615 256 8649 290
rect 8687 256 8721 290
rect 8759 256 8793 290
rect 8831 256 8865 290
rect 8903 256 8937 290
rect 9083 256 9117 290
rect 9155 256 9189 290
rect 9227 256 9261 290
rect 9299 256 9333 290
rect 9371 256 9405 290
rect 9443 256 9477 290
rect 9515 256 9549 290
rect 9587 256 9621 290
rect 9659 256 9693 290
rect 9731 256 9765 290
rect 9803 256 9837 290
rect 9983 256 10017 290
rect 10055 256 10089 290
rect 10127 256 10161 290
rect 10199 256 10233 290
rect 10271 256 10305 290
rect 10343 256 10377 290
rect 10415 256 10449 290
rect 10487 256 10521 290
rect 10559 256 10593 290
rect 10631 256 10665 290
rect 10703 256 10737 290
rect 10883 256 10917 290
rect 10955 256 10989 290
rect 11027 256 11061 290
rect 11099 256 11133 290
rect 11171 256 11205 290
rect 11243 256 11277 290
rect 11315 256 11349 290
rect 11387 256 11421 290
rect 11459 256 11493 290
rect 11531 256 11565 290
rect 11603 256 11637 290
rect 11783 256 11817 290
rect 11855 256 11889 290
rect 11927 256 11961 290
rect 11999 256 12033 290
rect 12071 256 12105 290
rect 12143 256 12177 290
rect 12215 256 12249 290
rect 12287 256 12321 290
rect 12359 256 12393 290
rect 12431 256 12465 290
rect 12503 256 12537 290
<< locali >>
rect 67 256 83 290
rect 117 256 155 290
rect 189 256 227 290
rect 261 256 299 290
rect 333 256 371 290
rect 405 256 443 290
rect 477 256 515 290
rect 549 256 587 290
rect 621 256 659 290
rect 693 256 731 290
rect 765 256 803 290
rect 837 256 853 290
rect 967 256 983 290
rect 1017 256 1055 290
rect 1089 256 1127 290
rect 1161 256 1199 290
rect 1233 256 1271 290
rect 1305 256 1343 290
rect 1377 256 1415 290
rect 1449 256 1487 290
rect 1521 256 1559 290
rect 1593 256 1631 290
rect 1665 256 1703 290
rect 1737 256 1753 290
rect 1867 256 1883 290
rect 1917 256 1955 290
rect 1989 256 2027 290
rect 2061 256 2099 290
rect 2133 256 2171 290
rect 2205 256 2243 290
rect 2277 256 2315 290
rect 2349 256 2387 290
rect 2421 256 2459 290
rect 2493 256 2531 290
rect 2565 256 2603 290
rect 2637 256 2653 290
rect 2767 256 2783 290
rect 2817 256 2855 290
rect 2889 256 2927 290
rect 2961 256 2999 290
rect 3033 256 3071 290
rect 3105 256 3143 290
rect 3177 256 3215 290
rect 3249 256 3287 290
rect 3321 256 3359 290
rect 3393 256 3431 290
rect 3465 256 3503 290
rect 3537 256 3553 290
rect 3667 256 3683 290
rect 3717 256 3755 290
rect 3789 256 3827 290
rect 3861 256 3899 290
rect 3933 256 3971 290
rect 4005 256 4043 290
rect 4077 256 4115 290
rect 4149 256 4187 290
rect 4221 256 4259 290
rect 4293 256 4331 290
rect 4365 256 4403 290
rect 4437 256 4453 290
rect 4567 256 4583 290
rect 4617 256 4655 290
rect 4689 256 4727 290
rect 4761 256 4799 290
rect 4833 256 4871 290
rect 4905 256 4943 290
rect 4977 256 5015 290
rect 5049 256 5087 290
rect 5121 256 5159 290
rect 5193 256 5231 290
rect 5265 256 5303 290
rect 5337 256 5353 290
rect 5467 256 5483 290
rect 5517 256 5555 290
rect 5589 256 5627 290
rect 5661 256 5699 290
rect 5733 256 5771 290
rect 5805 256 5843 290
rect 5877 256 5915 290
rect 5949 256 5987 290
rect 6021 256 6059 290
rect 6093 256 6131 290
rect 6165 256 6203 290
rect 6237 256 6253 290
rect 6367 256 6383 290
rect 6417 256 6455 290
rect 6489 256 6527 290
rect 6561 256 6599 290
rect 6633 256 6671 290
rect 6705 256 6743 290
rect 6777 256 6815 290
rect 6849 256 6887 290
rect 6921 256 6959 290
rect 6993 256 7031 290
rect 7065 256 7103 290
rect 7137 256 7153 290
rect 7267 256 7283 290
rect 7317 256 7355 290
rect 7389 256 7427 290
rect 7461 256 7499 290
rect 7533 256 7571 290
rect 7605 256 7643 290
rect 7677 256 7715 290
rect 7749 256 7787 290
rect 7821 256 7859 290
rect 7893 256 7931 290
rect 7965 256 8003 290
rect 8037 256 8053 290
rect 8167 256 8183 290
rect 8217 256 8255 290
rect 8289 256 8327 290
rect 8361 256 8399 290
rect 8433 256 8471 290
rect 8505 256 8543 290
rect 8577 256 8615 290
rect 8649 256 8687 290
rect 8721 256 8759 290
rect 8793 256 8831 290
rect 8865 256 8903 290
rect 8937 256 8953 290
rect 9067 256 9083 290
rect 9117 256 9155 290
rect 9189 256 9227 290
rect 9261 256 9299 290
rect 9333 256 9371 290
rect 9405 256 9443 290
rect 9477 256 9515 290
rect 9549 256 9587 290
rect 9621 256 9659 290
rect 9693 256 9731 290
rect 9765 256 9803 290
rect 9837 256 9853 290
rect 9967 256 9983 290
rect 10017 256 10055 290
rect 10089 256 10127 290
rect 10161 256 10199 290
rect 10233 256 10271 290
rect 10305 256 10343 290
rect 10377 256 10415 290
rect 10449 256 10487 290
rect 10521 256 10559 290
rect 10593 256 10631 290
rect 10665 256 10703 290
rect 10737 256 10753 290
rect 10867 256 10883 290
rect 10917 256 10955 290
rect 10989 256 11027 290
rect 11061 256 11099 290
rect 11133 256 11171 290
rect 11205 256 11243 290
rect 11277 256 11315 290
rect 11349 256 11387 290
rect 11421 256 11459 290
rect 11493 256 11531 290
rect 11565 256 11603 290
rect 11637 256 11653 290
rect 11767 256 11783 290
rect 11817 256 11855 290
rect 11889 256 11927 290
rect 11961 256 11999 290
rect 12033 256 12071 290
rect 12105 256 12143 290
rect 12177 256 12215 290
rect 12249 256 12287 290
rect 12321 256 12359 290
rect 12393 256 12431 290
rect 12465 256 12503 290
rect 12537 256 12553 290
rect 13 153 47 169
rect 13 81 47 119
rect 13 31 47 47
rect 893 153 927 169
rect 893 81 927 119
rect 893 31 927 47
rect 1793 153 1827 169
rect 1793 81 1827 119
rect 1793 31 1827 47
rect 2693 153 2727 169
rect 2693 81 2727 119
rect 2693 31 2727 47
rect 3593 153 3627 169
rect 3593 81 3627 119
rect 3593 31 3627 47
rect 4493 153 4527 169
rect 4493 81 4527 119
rect 4493 31 4527 47
rect 5393 153 5427 169
rect 5393 81 5427 119
rect 5393 31 5427 47
rect 6293 153 6327 169
rect 6293 81 6327 119
rect 6293 31 6327 47
rect 7193 153 7227 169
rect 7193 81 7227 119
rect 7193 31 7227 47
rect 8093 153 8127 169
rect 8093 81 8127 119
rect 8093 31 8127 47
rect 8993 153 9027 169
rect 8993 81 9027 119
rect 8993 31 9027 47
rect 9893 153 9927 169
rect 9893 81 9927 119
rect 9893 31 9927 47
rect 10793 153 10827 169
rect 10793 81 10827 119
rect 10793 31 10827 47
rect 11693 153 11727 169
rect 11693 81 11727 119
rect 11693 31 11727 47
rect 12573 153 12607 169
rect 12573 81 12607 119
rect 12573 31 12607 47
<< viali >>
rect 83 256 117 290
rect 155 256 189 290
rect 227 256 261 290
rect 299 256 333 290
rect 371 256 405 290
rect 443 256 477 290
rect 515 256 549 290
rect 587 256 621 290
rect 659 256 693 290
rect 731 256 765 290
rect 803 256 837 290
rect 983 256 1017 290
rect 1055 256 1089 290
rect 1127 256 1161 290
rect 1199 256 1233 290
rect 1271 256 1305 290
rect 1343 256 1377 290
rect 1415 256 1449 290
rect 1487 256 1521 290
rect 1559 256 1593 290
rect 1631 256 1665 290
rect 1703 256 1737 290
rect 1883 256 1917 290
rect 1955 256 1989 290
rect 2027 256 2061 290
rect 2099 256 2133 290
rect 2171 256 2205 290
rect 2243 256 2277 290
rect 2315 256 2349 290
rect 2387 256 2421 290
rect 2459 256 2493 290
rect 2531 256 2565 290
rect 2603 256 2637 290
rect 2783 256 2817 290
rect 2855 256 2889 290
rect 2927 256 2961 290
rect 2999 256 3033 290
rect 3071 256 3105 290
rect 3143 256 3177 290
rect 3215 256 3249 290
rect 3287 256 3321 290
rect 3359 256 3393 290
rect 3431 256 3465 290
rect 3503 256 3537 290
rect 3683 256 3717 290
rect 3755 256 3789 290
rect 3827 256 3861 290
rect 3899 256 3933 290
rect 3971 256 4005 290
rect 4043 256 4077 290
rect 4115 256 4149 290
rect 4187 256 4221 290
rect 4259 256 4293 290
rect 4331 256 4365 290
rect 4403 256 4437 290
rect 4583 256 4617 290
rect 4655 256 4689 290
rect 4727 256 4761 290
rect 4799 256 4833 290
rect 4871 256 4905 290
rect 4943 256 4977 290
rect 5015 256 5049 290
rect 5087 256 5121 290
rect 5159 256 5193 290
rect 5231 256 5265 290
rect 5303 256 5337 290
rect 5483 256 5517 290
rect 5555 256 5589 290
rect 5627 256 5661 290
rect 5699 256 5733 290
rect 5771 256 5805 290
rect 5843 256 5877 290
rect 5915 256 5949 290
rect 5987 256 6021 290
rect 6059 256 6093 290
rect 6131 256 6165 290
rect 6203 256 6237 290
rect 6383 256 6417 290
rect 6455 256 6489 290
rect 6527 256 6561 290
rect 6599 256 6633 290
rect 6671 256 6705 290
rect 6743 256 6777 290
rect 6815 256 6849 290
rect 6887 256 6921 290
rect 6959 256 6993 290
rect 7031 256 7065 290
rect 7103 256 7137 290
rect 7283 256 7317 290
rect 7355 256 7389 290
rect 7427 256 7461 290
rect 7499 256 7533 290
rect 7571 256 7605 290
rect 7643 256 7677 290
rect 7715 256 7749 290
rect 7787 256 7821 290
rect 7859 256 7893 290
rect 7931 256 7965 290
rect 8003 256 8037 290
rect 8183 256 8217 290
rect 8255 256 8289 290
rect 8327 256 8361 290
rect 8399 256 8433 290
rect 8471 256 8505 290
rect 8543 256 8577 290
rect 8615 256 8649 290
rect 8687 256 8721 290
rect 8759 256 8793 290
rect 8831 256 8865 290
rect 8903 256 8937 290
rect 9083 256 9117 290
rect 9155 256 9189 290
rect 9227 256 9261 290
rect 9299 256 9333 290
rect 9371 256 9405 290
rect 9443 256 9477 290
rect 9515 256 9549 290
rect 9587 256 9621 290
rect 9659 256 9693 290
rect 9731 256 9765 290
rect 9803 256 9837 290
rect 9983 256 10017 290
rect 10055 256 10089 290
rect 10127 256 10161 290
rect 10199 256 10233 290
rect 10271 256 10305 290
rect 10343 256 10377 290
rect 10415 256 10449 290
rect 10487 256 10521 290
rect 10559 256 10593 290
rect 10631 256 10665 290
rect 10703 256 10737 290
rect 10883 256 10917 290
rect 10955 256 10989 290
rect 11027 256 11061 290
rect 11099 256 11133 290
rect 11171 256 11205 290
rect 11243 256 11277 290
rect 11315 256 11349 290
rect 11387 256 11421 290
rect 11459 256 11493 290
rect 11531 256 11565 290
rect 11603 256 11637 290
rect 11783 256 11817 290
rect 11855 256 11889 290
rect 11927 256 11961 290
rect 11999 256 12033 290
rect 12071 256 12105 290
rect 12143 256 12177 290
rect 12215 256 12249 290
rect 12287 256 12321 290
rect 12359 256 12393 290
rect 12431 256 12465 290
rect 12503 256 12537 290
rect 13 119 47 153
rect 13 47 47 81
rect 893 119 927 153
rect 893 47 927 81
rect 1793 119 1827 153
rect 1793 47 1827 81
rect 2693 119 2727 153
rect 2693 47 2727 81
rect 3593 119 3627 153
rect 3593 47 3627 81
rect 4493 119 4527 153
rect 4493 47 4527 81
rect 5393 119 5427 153
rect 5393 47 5427 81
rect 6293 119 6327 153
rect 6293 47 6327 81
rect 7193 119 7227 153
rect 7193 47 7227 81
rect 8093 119 8127 153
rect 8093 47 8127 81
rect 8993 119 9027 153
rect 8993 47 9027 81
rect 9893 119 9927 153
rect 9893 47 9927 81
rect 10793 119 10827 153
rect 10793 47 10827 81
rect 11693 119 11727 153
rect 11693 47 11727 81
rect 12573 119 12607 153
rect 12573 47 12607 81
<< metal1 >>
rect 71 290 849 296
rect 71 256 83 290
rect 117 256 155 290
rect 189 256 227 290
rect 261 256 299 290
rect 333 256 371 290
rect 405 256 443 290
rect 477 256 515 290
rect 549 256 587 290
rect 621 256 659 290
rect 693 256 731 290
rect 765 256 803 290
rect 837 256 849 290
rect 71 250 849 256
rect 971 290 1749 296
rect 971 256 983 290
rect 1017 256 1055 290
rect 1089 256 1127 290
rect 1161 256 1199 290
rect 1233 256 1271 290
rect 1305 256 1343 290
rect 1377 256 1415 290
rect 1449 256 1487 290
rect 1521 256 1559 290
rect 1593 256 1631 290
rect 1665 256 1703 290
rect 1737 256 1749 290
rect 971 250 1749 256
rect 1871 290 2649 296
rect 1871 256 1883 290
rect 1917 256 1955 290
rect 1989 256 2027 290
rect 2061 256 2099 290
rect 2133 256 2171 290
rect 2205 256 2243 290
rect 2277 256 2315 290
rect 2349 256 2387 290
rect 2421 256 2459 290
rect 2493 256 2531 290
rect 2565 256 2603 290
rect 2637 256 2649 290
rect 1871 250 2649 256
rect 2771 290 3549 296
rect 2771 256 2783 290
rect 2817 256 2855 290
rect 2889 256 2927 290
rect 2961 256 2999 290
rect 3033 256 3071 290
rect 3105 256 3143 290
rect 3177 256 3215 290
rect 3249 256 3287 290
rect 3321 256 3359 290
rect 3393 256 3431 290
rect 3465 256 3503 290
rect 3537 256 3549 290
rect 2771 250 3549 256
rect 3671 290 4449 296
rect 3671 256 3683 290
rect 3717 256 3755 290
rect 3789 256 3827 290
rect 3861 256 3899 290
rect 3933 256 3971 290
rect 4005 256 4043 290
rect 4077 256 4115 290
rect 4149 256 4187 290
rect 4221 256 4259 290
rect 4293 256 4331 290
rect 4365 256 4403 290
rect 4437 256 4449 290
rect 3671 250 4449 256
rect 4571 290 5349 296
rect 4571 256 4583 290
rect 4617 256 4655 290
rect 4689 256 4727 290
rect 4761 256 4799 290
rect 4833 256 4871 290
rect 4905 256 4943 290
rect 4977 256 5015 290
rect 5049 256 5087 290
rect 5121 256 5159 290
rect 5193 256 5231 290
rect 5265 256 5303 290
rect 5337 256 5349 290
rect 4571 250 5349 256
rect 5471 290 6249 296
rect 5471 256 5483 290
rect 5517 256 5555 290
rect 5589 256 5627 290
rect 5661 256 5699 290
rect 5733 256 5771 290
rect 5805 256 5843 290
rect 5877 256 5915 290
rect 5949 256 5987 290
rect 6021 256 6059 290
rect 6093 256 6131 290
rect 6165 256 6203 290
rect 6237 256 6249 290
rect 5471 250 6249 256
rect 6371 290 7149 296
rect 6371 256 6383 290
rect 6417 256 6455 290
rect 6489 256 6527 290
rect 6561 256 6599 290
rect 6633 256 6671 290
rect 6705 256 6743 290
rect 6777 256 6815 290
rect 6849 256 6887 290
rect 6921 256 6959 290
rect 6993 256 7031 290
rect 7065 256 7103 290
rect 7137 256 7149 290
rect 6371 250 7149 256
rect 7271 290 8049 296
rect 7271 256 7283 290
rect 7317 256 7355 290
rect 7389 256 7427 290
rect 7461 256 7499 290
rect 7533 256 7571 290
rect 7605 256 7643 290
rect 7677 256 7715 290
rect 7749 256 7787 290
rect 7821 256 7859 290
rect 7893 256 7931 290
rect 7965 256 8003 290
rect 8037 256 8049 290
rect 7271 250 8049 256
rect 8171 290 8949 296
rect 8171 256 8183 290
rect 8217 256 8255 290
rect 8289 256 8327 290
rect 8361 256 8399 290
rect 8433 256 8471 290
rect 8505 256 8543 290
rect 8577 256 8615 290
rect 8649 256 8687 290
rect 8721 256 8759 290
rect 8793 256 8831 290
rect 8865 256 8903 290
rect 8937 256 8949 290
rect 8171 250 8949 256
rect 9071 290 9849 296
rect 9071 256 9083 290
rect 9117 256 9155 290
rect 9189 256 9227 290
rect 9261 256 9299 290
rect 9333 256 9371 290
rect 9405 256 9443 290
rect 9477 256 9515 290
rect 9549 256 9587 290
rect 9621 256 9659 290
rect 9693 256 9731 290
rect 9765 256 9803 290
rect 9837 256 9849 290
rect 9071 250 9849 256
rect 9971 290 10749 296
rect 9971 256 9983 290
rect 10017 256 10055 290
rect 10089 256 10127 290
rect 10161 256 10199 290
rect 10233 256 10271 290
rect 10305 256 10343 290
rect 10377 256 10415 290
rect 10449 256 10487 290
rect 10521 256 10559 290
rect 10593 256 10631 290
rect 10665 256 10703 290
rect 10737 256 10749 290
rect 9971 250 10749 256
rect 10871 290 11649 296
rect 10871 256 10883 290
rect 10917 256 10955 290
rect 10989 256 11027 290
rect 11061 256 11099 290
rect 11133 256 11171 290
rect 11205 256 11243 290
rect 11277 256 11315 290
rect 11349 256 11387 290
rect 11421 256 11459 290
rect 11493 256 11531 290
rect 11565 256 11603 290
rect 11637 256 11649 290
rect 10871 250 11649 256
rect 11771 290 12549 296
rect 11771 256 11783 290
rect 11817 256 11855 290
rect 11889 256 11927 290
rect 11961 256 11999 290
rect 12033 256 12071 290
rect 12105 256 12143 290
rect 12177 256 12215 290
rect 12249 256 12287 290
rect 12321 256 12359 290
rect 12393 256 12431 290
rect 12465 256 12503 290
rect 12537 256 12549 290
rect 11771 250 12549 256
rect 7 153 53 165
rect 7 119 13 153
rect 47 119 53 153
rect 7 81 53 119
rect 7 47 13 81
rect 47 47 53 81
rect 7 35 53 47
rect 887 153 933 165
rect 887 119 893 153
rect 927 119 933 153
rect 887 81 933 119
rect 887 47 893 81
rect 927 47 933 81
rect 887 35 933 47
rect 1787 153 1833 165
rect 1787 119 1793 153
rect 1827 119 1833 153
rect 1787 81 1833 119
rect 1787 47 1793 81
rect 1827 47 1833 81
rect 1787 35 1833 47
rect 2687 153 2733 165
rect 2687 119 2693 153
rect 2727 119 2733 153
rect 2687 81 2733 119
rect 2687 47 2693 81
rect 2727 47 2733 81
rect 2687 35 2733 47
rect 3587 153 3633 165
rect 3587 119 3593 153
rect 3627 119 3633 153
rect 3587 81 3633 119
rect 3587 47 3593 81
rect 3627 47 3633 81
rect 3587 35 3633 47
rect 4487 153 4533 165
rect 4487 119 4493 153
rect 4527 119 4533 153
rect 4487 81 4533 119
rect 4487 47 4493 81
rect 4527 47 4533 81
rect 4487 35 4533 47
rect 5387 153 5433 165
rect 5387 119 5393 153
rect 5427 119 5433 153
rect 5387 81 5433 119
rect 5387 47 5393 81
rect 5427 47 5433 81
rect 5387 35 5433 47
rect 6287 153 6333 165
rect 6287 119 6293 153
rect 6327 119 6333 153
rect 6287 81 6333 119
rect 6287 47 6293 81
rect 6327 47 6333 81
rect 6287 35 6333 47
rect 7187 153 7233 165
rect 7187 119 7193 153
rect 7227 119 7233 153
rect 7187 81 7233 119
rect 7187 47 7193 81
rect 7227 47 7233 81
rect 7187 35 7233 47
rect 8087 153 8133 165
rect 8087 119 8093 153
rect 8127 119 8133 153
rect 8087 81 8133 119
rect 8087 47 8093 81
rect 8127 47 8133 81
rect 8087 35 8133 47
rect 8987 153 9033 165
rect 8987 119 8993 153
rect 9027 119 9033 153
rect 8987 81 9033 119
rect 8987 47 8993 81
rect 9027 47 9033 81
rect 8987 35 9033 47
rect 9887 153 9933 165
rect 9887 119 9893 153
rect 9927 119 9933 153
rect 9887 81 9933 119
rect 9887 47 9893 81
rect 9927 47 9933 81
rect 9887 35 9933 47
rect 10787 153 10833 165
rect 10787 119 10793 153
rect 10827 119 10833 153
rect 10787 81 10833 119
rect 10787 47 10793 81
rect 10827 47 10833 81
rect 10787 35 10833 47
rect 11687 153 11733 165
rect 11687 119 11693 153
rect 11727 119 11733 153
rect 11687 81 11733 119
rect 11687 47 11693 81
rect 11727 47 11733 81
rect 11687 35 11733 47
rect 12567 153 12613 165
rect 12567 119 12573 153
rect 12607 119 12613 153
rect 12567 81 12613 119
rect 12567 47 12573 81
rect 12607 47 12613 81
rect 12567 35 12613 47
<< end >>
