magic
tech sky130A
magscale 1 2
timestamp 1693698878
<< nwell >>
rect -338 -6887 338 6887
<< mvpmos >>
rect -80 4590 80 6590
rect -80 2354 80 4354
rect -80 118 80 2118
rect -80 -2118 80 -118
rect -80 -4354 80 -2354
rect -80 -6590 80 -4590
<< mvpdiff >>
rect -138 6578 -80 6590
rect -138 4602 -126 6578
rect -92 4602 -80 6578
rect -138 4590 -80 4602
rect 80 6578 138 6590
rect 80 4602 92 6578
rect 126 4602 138 6578
rect 80 4590 138 4602
rect -138 4342 -80 4354
rect -138 2366 -126 4342
rect -92 2366 -80 4342
rect -138 2354 -80 2366
rect 80 4342 138 4354
rect 80 2366 92 4342
rect 126 2366 138 4342
rect 80 2354 138 2366
rect -138 2106 -80 2118
rect -138 130 -126 2106
rect -92 130 -80 2106
rect -138 118 -80 130
rect 80 2106 138 2118
rect 80 130 92 2106
rect 126 130 138 2106
rect 80 118 138 130
rect -138 -130 -80 -118
rect -138 -2106 -126 -130
rect -92 -2106 -80 -130
rect -138 -2118 -80 -2106
rect 80 -130 138 -118
rect 80 -2106 92 -130
rect 126 -2106 138 -130
rect 80 -2118 138 -2106
rect -138 -2366 -80 -2354
rect -138 -4342 -126 -2366
rect -92 -4342 -80 -2366
rect -138 -4354 -80 -4342
rect 80 -2366 138 -2354
rect 80 -4342 92 -2366
rect 126 -4342 138 -2366
rect 80 -4354 138 -4342
rect -138 -4602 -80 -4590
rect -138 -6578 -126 -4602
rect -92 -6578 -80 -4602
rect -138 -6590 -80 -6578
rect 80 -4602 138 -4590
rect 80 -6578 92 -4602
rect 126 -6578 138 -4602
rect 80 -6590 138 -6578
<< mvpdiffc >>
rect -126 4602 -92 6578
rect 92 4602 126 6578
rect -126 2366 -92 4342
rect 92 2366 126 4342
rect -126 130 -92 2106
rect 92 130 126 2106
rect -126 -2106 -92 -130
rect 92 -2106 126 -130
rect -126 -4342 -92 -2366
rect 92 -4342 126 -2366
rect -126 -6578 -92 -4602
rect 92 -6578 126 -4602
<< mvnsubdiff >>
rect -272 6809 272 6821
rect -272 6775 -164 6809
rect 164 6775 272 6809
rect -272 6763 272 6775
rect -272 6713 -214 6763
rect -272 -6713 -260 6713
rect -226 -6713 -214 6713
rect 214 6713 272 6763
rect -272 -6763 -214 -6713
rect 214 -6713 226 6713
rect 260 -6713 272 6713
rect 214 -6763 272 -6713
rect -272 -6775 272 -6763
rect -272 -6809 -164 -6775
rect 164 -6809 272 -6775
rect -272 -6821 272 -6809
<< mvnsubdiffcont >>
rect -164 6775 164 6809
rect -260 -6713 -226 6713
rect 226 -6713 260 6713
rect -164 -6809 164 -6775
<< poly >>
rect -80 6671 80 6687
rect -80 6637 -64 6671
rect 64 6637 80 6671
rect -80 6590 80 6637
rect -80 4543 80 4590
rect -80 4509 -64 4543
rect 64 4509 80 4543
rect -80 4493 80 4509
rect -80 4435 80 4451
rect -80 4401 -64 4435
rect 64 4401 80 4435
rect -80 4354 80 4401
rect -80 2307 80 2354
rect -80 2273 -64 2307
rect 64 2273 80 2307
rect -80 2257 80 2273
rect -80 2199 80 2215
rect -80 2165 -64 2199
rect 64 2165 80 2199
rect -80 2118 80 2165
rect -80 71 80 118
rect -80 37 -64 71
rect 64 37 80 71
rect -80 21 80 37
rect -80 -37 80 -21
rect -80 -71 -64 -37
rect 64 -71 80 -37
rect -80 -118 80 -71
rect -80 -2165 80 -2118
rect -80 -2199 -64 -2165
rect 64 -2199 80 -2165
rect -80 -2215 80 -2199
rect -80 -2273 80 -2257
rect -80 -2307 -64 -2273
rect 64 -2307 80 -2273
rect -80 -2354 80 -2307
rect -80 -4401 80 -4354
rect -80 -4435 -64 -4401
rect 64 -4435 80 -4401
rect -80 -4451 80 -4435
rect -80 -4509 80 -4493
rect -80 -4543 -64 -4509
rect 64 -4543 80 -4509
rect -80 -4590 80 -4543
rect -80 -6637 80 -6590
rect -80 -6671 -64 -6637
rect 64 -6671 80 -6637
rect -80 -6687 80 -6671
<< polycont >>
rect -64 6637 64 6671
rect -64 4509 64 4543
rect -64 4401 64 4435
rect -64 2273 64 2307
rect -64 2165 64 2199
rect -64 37 64 71
rect -64 -71 64 -37
rect -64 -2199 64 -2165
rect -64 -2307 64 -2273
rect -64 -4435 64 -4401
rect -64 -4543 64 -4509
rect -64 -6671 64 -6637
<< locali >>
rect -260 6775 -164 6809
rect 164 6775 260 6809
rect -260 6713 -226 6775
rect 226 6713 260 6775
rect -80 6637 -64 6671
rect 64 6637 80 6671
rect -126 6578 -92 6594
rect -126 4586 -92 4602
rect 92 6578 126 6594
rect 92 4586 126 4602
rect -80 4509 -64 4543
rect 64 4509 80 4543
rect -80 4401 -64 4435
rect 64 4401 80 4435
rect -126 4342 -92 4358
rect -126 2350 -92 2366
rect 92 4342 126 4358
rect 92 2350 126 2366
rect -80 2273 -64 2307
rect 64 2273 80 2307
rect -80 2165 -64 2199
rect 64 2165 80 2199
rect -126 2106 -92 2122
rect -126 114 -92 130
rect 92 2106 126 2122
rect 92 114 126 130
rect -80 37 -64 71
rect 64 37 80 71
rect -80 -71 -64 -37
rect 64 -71 80 -37
rect -126 -130 -92 -114
rect -126 -2122 -92 -2106
rect 92 -130 126 -114
rect 92 -2122 126 -2106
rect -80 -2199 -64 -2165
rect 64 -2199 80 -2165
rect -80 -2307 -64 -2273
rect 64 -2307 80 -2273
rect -126 -2366 -92 -2350
rect -126 -4358 -92 -4342
rect 92 -2366 126 -2350
rect 92 -4358 126 -4342
rect -80 -4435 -64 -4401
rect 64 -4435 80 -4401
rect -80 -4543 -64 -4509
rect 64 -4543 80 -4509
rect -126 -4602 -92 -4586
rect -126 -6594 -92 -6578
rect 92 -4602 126 -4586
rect 92 -6594 126 -6578
rect -80 -6671 -64 -6637
rect 64 -6671 80 -6637
rect -260 -6775 -226 -6713
rect 226 -6775 260 -6713
rect -260 -6809 -164 -6775
rect 164 -6809 260 -6775
<< viali >>
rect -64 6637 64 6671
rect -126 4602 -92 6578
rect 92 4602 126 6578
rect -64 4509 64 4543
rect -64 4401 64 4435
rect -126 2366 -92 4342
rect 92 2366 126 4342
rect -64 2273 64 2307
rect -64 2165 64 2199
rect -126 130 -92 2106
rect 92 130 126 2106
rect -64 37 64 71
rect -64 -71 64 -37
rect -126 -2106 -92 -130
rect 92 -2106 126 -130
rect -64 -2199 64 -2165
rect -64 -2307 64 -2273
rect -126 -4342 -92 -2366
rect 92 -4342 126 -2366
rect -64 -4435 64 -4401
rect -64 -4543 64 -4509
rect -126 -6578 -92 -4602
rect 92 -6578 126 -4602
rect -64 -6671 64 -6637
<< metal1 >>
rect -76 6671 76 6677
rect -76 6637 -64 6671
rect 64 6637 76 6671
rect -76 6631 76 6637
rect -132 6578 -86 6590
rect -132 4602 -126 6578
rect -92 4602 -86 6578
rect -132 4590 -86 4602
rect 86 6578 132 6590
rect 86 4602 92 6578
rect 126 4602 132 6578
rect 86 4590 132 4602
rect -76 4543 76 4549
rect -76 4509 -64 4543
rect 64 4509 76 4543
rect -76 4503 76 4509
rect -76 4435 76 4441
rect -76 4401 -64 4435
rect 64 4401 76 4435
rect -76 4395 76 4401
rect -132 4342 -86 4354
rect -132 2366 -126 4342
rect -92 2366 -86 4342
rect -132 2354 -86 2366
rect 86 4342 132 4354
rect 86 2366 92 4342
rect 126 2366 132 4342
rect 86 2354 132 2366
rect -76 2307 76 2313
rect -76 2273 -64 2307
rect 64 2273 76 2307
rect -76 2267 76 2273
rect -76 2199 76 2205
rect -76 2165 -64 2199
rect 64 2165 76 2199
rect -76 2159 76 2165
rect -132 2106 -86 2118
rect -132 130 -126 2106
rect -92 130 -86 2106
rect -132 118 -86 130
rect 86 2106 132 2118
rect 86 130 92 2106
rect 126 130 132 2106
rect 86 118 132 130
rect -76 71 76 77
rect -76 37 -64 71
rect 64 37 76 71
rect -76 31 76 37
rect -76 -37 76 -31
rect -76 -71 -64 -37
rect 64 -71 76 -37
rect -76 -77 76 -71
rect -132 -130 -86 -118
rect -132 -2106 -126 -130
rect -92 -2106 -86 -130
rect -132 -2118 -86 -2106
rect 86 -130 132 -118
rect 86 -2106 92 -130
rect 126 -2106 132 -130
rect 86 -2118 132 -2106
rect -76 -2165 76 -2159
rect -76 -2199 -64 -2165
rect 64 -2199 76 -2165
rect -76 -2205 76 -2199
rect -76 -2273 76 -2267
rect -76 -2307 -64 -2273
rect 64 -2307 76 -2273
rect -76 -2313 76 -2307
rect -132 -2366 -86 -2354
rect -132 -4342 -126 -2366
rect -92 -4342 -86 -2366
rect -132 -4354 -86 -4342
rect 86 -2366 132 -2354
rect 86 -4342 92 -2366
rect 126 -4342 132 -2366
rect 86 -4354 132 -4342
rect -76 -4401 76 -4395
rect -76 -4435 -64 -4401
rect 64 -4435 76 -4401
rect -76 -4441 76 -4435
rect -76 -4509 76 -4503
rect -76 -4543 -64 -4509
rect 64 -4543 76 -4509
rect -76 -4549 76 -4543
rect -132 -4602 -86 -4590
rect -132 -6578 -126 -4602
rect -92 -6578 -86 -4602
rect -132 -6590 -86 -6578
rect 86 -4602 132 -4590
rect 86 -6578 92 -4602
rect 126 -6578 132 -4602
rect 86 -6590 132 -6578
rect -76 -6637 76 -6631
rect -76 -6671 -64 -6637
rect 64 -6671 76 -6637
rect -76 -6677 76 -6671
<< properties >>
string FIXED_BBOX -243 -6792 243 6792
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 10 l 0.8 m 6 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
