magic
tech sky130A
magscale 1 2
timestamp 1740486730
<< xpolycontact >>
rect -35 164 35 596
rect -35 -596 35 -164
<< ppolyres >>
rect -35 -164 35 164
<< viali >>
rect -19 181 19 578
rect -19 -578 19 -181
<< metal1 >>
rect -25 578 25 590
rect -25 181 -19 578
rect 19 181 25 578
rect -25 169 25 181
rect -25 -181 25 -169
rect -25 -578 -19 -181
rect 19 -578 25 -181
rect -25 -590 25 -578
<< properties >>
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 1.8 m 1 nx 1 wmin 0.350 lmin 0.50 class resistor rho 319.8 val 2.757k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
