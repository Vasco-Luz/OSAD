magic
tech sky130A
magscale 1 2
timestamp 1740348852
<< error_p >>
rect -1091 -130 1091 202
rect -1061 -164 1061 -130
<< nwell >>
rect -1061 -164 1061 198
<< mvpmos >>
rect -967 -64 -527 136
rect -469 -64 -29 136
rect 29 -64 469 136
rect 527 -64 967 136
<< mvpdiff >>
rect -1025 124 -967 136
rect -1025 -52 -1013 124
rect -979 -52 -967 124
rect -1025 -64 -967 -52
rect -527 124 -469 136
rect -527 -52 -515 124
rect -481 -52 -469 124
rect -527 -64 -469 -52
rect -29 124 29 136
rect -29 -52 -17 124
rect 17 -52 29 124
rect -29 -64 29 -52
rect 469 124 527 136
rect 469 -52 481 124
rect 515 -52 527 124
rect 469 -64 527 -52
rect 967 124 1025 136
rect 967 -52 979 124
rect 1013 -52 1025 124
rect 967 -64 1025 -52
<< mvpdiffc >>
rect -1013 -52 -979 124
rect -515 -52 -481 124
rect -17 -52 17 124
rect 481 -52 515 124
rect 979 -52 1013 124
<< poly >>
rect -967 136 -527 162
rect -469 136 -29 162
rect 29 136 469 162
rect 527 136 967 162
rect -967 -111 -527 -64
rect -967 -128 -910 -111
rect -926 -145 -910 -128
rect -584 -128 -527 -111
rect -469 -111 -29 -64
rect -469 -128 -412 -111
rect -584 -145 -568 -128
rect -926 -161 -568 -145
rect -428 -145 -412 -128
rect -86 -128 -29 -111
rect 29 -111 469 -64
rect 29 -128 86 -111
rect -86 -145 -70 -128
rect -428 -161 -70 -145
rect 70 -145 86 -128
rect 412 -128 469 -111
rect 527 -111 967 -64
rect 527 -128 584 -111
rect 412 -145 428 -128
rect 70 -161 428 -145
rect 568 -145 584 -128
rect 910 -128 967 -111
rect 910 -145 926 -128
rect 568 -161 926 -145
<< polycont >>
rect -910 -145 -584 -111
rect -412 -145 -86 -111
rect 86 -145 412 -111
rect 584 -145 910 -111
<< locali >>
rect -1013 124 -979 140
rect -1013 -68 -979 -52
rect -515 124 -481 140
rect -515 -68 -481 -52
rect -17 124 17 140
rect -17 -68 17 -52
rect 481 124 515 140
rect 481 -68 515 -52
rect 979 124 1013 140
rect 979 -68 1013 -52
rect -927 -111 -567 -106
rect -927 -145 -910 -111
rect -584 -145 -567 -111
rect -927 -180 -567 -145
rect -429 -111 -69 -106
rect -429 -145 -412 -111
rect -86 -145 -69 -111
rect -429 -180 -69 -145
rect 69 -111 429 -106
rect 69 -145 86 -111
rect 412 -145 429 -111
rect 69 -180 429 -145
rect 567 -111 927 -106
rect 567 -145 584 -111
rect 910 -145 927 -111
rect 567 -180 927 -145
rect -1007 -239 1030 -180
rect -1007 -240 -567 -239
rect -429 -240 -69 -239
rect 69 -240 429 -239
rect 567 -240 995 -239
<< viali >>
rect -1013 -52 -979 124
rect -515 -52 -481 124
rect -17 -52 17 124
rect 481 -52 515 124
rect 979 -52 1013 124
rect -910 -145 -584 -111
rect -412 -145 -86 -111
rect 86 -145 412 -111
rect 584 -145 910 -111
<< metal1 >>
rect -1013 136 -979 218
rect -17 136 17 464
rect 979 136 1013 508
rect -1019 124 -973 136
rect -1019 -52 -1013 124
rect -979 -52 -973 124
rect -1019 -64 -973 -52
rect -521 124 -475 136
rect -521 -52 -515 124
rect -481 -52 -475 124
rect -521 -64 -475 -52
rect -23 124 23 136
rect -23 -52 -17 124
rect 17 -52 23 124
rect -23 -64 23 -52
rect 475 124 521 136
rect 475 -52 481 124
rect 515 -52 521 124
rect 475 -64 521 -52
rect 973 124 1019 136
rect 973 -52 979 124
rect 1013 -52 1019 124
rect 973 -64 1019 -52
rect -1013 -102 -979 -64
rect -922 -111 -572 -105
rect -922 -145 -910 -111
rect -584 -145 -572 -111
rect -922 -151 -572 -145
rect -515 -384 -481 -64
rect -424 -111 -74 -105
rect -424 -145 -412 -111
rect -86 -145 -74 -111
rect -424 -151 -74 -145
rect 74 -111 424 -105
rect 74 -145 86 -111
rect 412 -145 424 -111
rect 74 -151 424 -145
rect 481 -394 515 -64
rect 572 -111 922 -105
rect 572 -145 584 -111
rect 910 -145 922 -111
rect 572 -151 922 -145
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1 l 2.2 m 1 nf 4 diffcov 100 polycov 80 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 80 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
