magic
tech sky130A
magscale 1 2
timestamp 1740397409
<< error_p >>
rect -378 -131 -320 69
rect 320 -131 378 69
<< mvnmos >>
rect -320 -131 320 69
<< mvndiff >>
rect -378 57 -320 69
rect -378 -119 -366 57
rect -332 -119 -320 57
rect -378 -131 -320 -119
rect 320 57 378 69
rect 320 -119 332 57
rect 366 -119 378 57
rect 320 -131 378 -119
<< mvndiffc >>
rect -366 -119 -332 57
rect 332 -119 366 57
<< poly >>
rect -259 141 259 157
rect -259 124 -243 141
rect -320 107 -243 124
rect 243 124 259 141
rect 243 107 320 124
rect -320 69 320 107
rect -320 -157 320 -131
<< polycont >>
rect -243 107 243 141
<< locali >>
rect -259 107 -243 141
rect 243 107 259 141
rect -366 57 -332 73
rect -366 -135 -332 -119
rect 332 57 366 73
rect 332 -135 366 -119
<< viali >>
rect -243 107 243 141
rect -366 -119 -332 57
rect 332 -119 366 57
<< metal1 >>
rect -366 141 255 147
rect -366 107 -243 141
rect 243 107 255 141
rect -366 101 255 107
rect -366 69 -332 101
rect -372 57 -326 69
rect -372 -119 -366 57
rect -332 -119 -326 57
rect -372 -131 -326 -119
rect 326 57 372 69
rect 326 -119 332 57
rect 366 -119 372 57
rect 326 -131 372 -119
<< labels >>
flabel mvnmos -96 -65 14 11 0 FreeSans 1600 0 0 0 D
flabel mvnmos -88 -67 22 9 0 FreeSans 1600 0 0 0 D
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 1 l 3.2 m 1 nf 1 diffcov 100 polycov 80 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 80 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
