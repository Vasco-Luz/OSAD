magic
tech sky130A
magscale 1 2
timestamp 1693698878
<< nwell >>
rect -1537 -662 1537 662
<< mvpmos >>
rect -1279 -436 -1119 364
rect -1061 -436 -901 364
rect -843 -436 -683 364
rect -625 -436 -465 364
rect -407 -436 -247 364
rect -189 -436 -29 364
rect 29 -436 189 364
rect 247 -436 407 364
rect 465 -436 625 364
rect 683 -436 843 364
rect 901 -436 1061 364
rect 1119 -436 1279 364
<< mvpdiff >>
rect -1337 352 -1279 364
rect -1337 -424 -1325 352
rect -1291 -424 -1279 352
rect -1337 -436 -1279 -424
rect -1119 352 -1061 364
rect -1119 -424 -1107 352
rect -1073 -424 -1061 352
rect -1119 -436 -1061 -424
rect -901 352 -843 364
rect -901 -424 -889 352
rect -855 -424 -843 352
rect -901 -436 -843 -424
rect -683 352 -625 364
rect -683 -424 -671 352
rect -637 -424 -625 352
rect -683 -436 -625 -424
rect -465 352 -407 364
rect -465 -424 -453 352
rect -419 -424 -407 352
rect -465 -436 -407 -424
rect -247 352 -189 364
rect -247 -424 -235 352
rect -201 -424 -189 352
rect -247 -436 -189 -424
rect -29 352 29 364
rect -29 -424 -17 352
rect 17 -424 29 352
rect -29 -436 29 -424
rect 189 352 247 364
rect 189 -424 201 352
rect 235 -424 247 352
rect 189 -436 247 -424
rect 407 352 465 364
rect 407 -424 419 352
rect 453 -424 465 352
rect 407 -436 465 -424
rect 625 352 683 364
rect 625 -424 637 352
rect 671 -424 683 352
rect 625 -436 683 -424
rect 843 352 901 364
rect 843 -424 855 352
rect 889 -424 901 352
rect 843 -436 901 -424
rect 1061 352 1119 364
rect 1061 -424 1073 352
rect 1107 -424 1119 352
rect 1061 -436 1119 -424
rect 1279 352 1337 364
rect 1279 -424 1291 352
rect 1325 -424 1337 352
rect 1279 -436 1337 -424
<< mvpdiffc >>
rect -1325 -424 -1291 352
rect -1107 -424 -1073 352
rect -889 -424 -855 352
rect -671 -424 -637 352
rect -453 -424 -419 352
rect -235 -424 -201 352
rect -17 -424 17 352
rect 201 -424 235 352
rect 419 -424 453 352
rect 637 -424 671 352
rect 855 -424 889 352
rect 1073 -424 1107 352
rect 1291 -424 1325 352
<< mvnsubdiff >>
rect -1471 584 1471 596
rect -1471 550 -1363 584
rect 1363 550 1471 584
rect -1471 538 1471 550
rect -1471 488 -1413 538
rect -1471 -488 -1459 488
rect -1425 -488 -1413 488
rect 1413 488 1471 538
rect -1471 -538 -1413 -488
rect 1413 -488 1425 488
rect 1459 -488 1471 488
rect 1413 -538 1471 -488
rect -1471 -550 1471 -538
rect -1471 -584 -1363 -550
rect 1363 -584 1471 -550
rect -1471 -596 1471 -584
<< mvnsubdiffcont >>
rect -1363 550 1363 584
rect -1459 -488 -1425 488
rect 1425 -488 1459 488
rect -1363 -584 1363 -550
<< poly >>
rect -1279 445 -1119 461
rect -1279 411 -1263 445
rect -1135 411 -1119 445
rect -1279 364 -1119 411
rect -1061 445 -901 461
rect -1061 411 -1045 445
rect -917 411 -901 445
rect -1061 364 -901 411
rect -843 445 -683 461
rect -843 411 -827 445
rect -699 411 -683 445
rect -843 364 -683 411
rect -625 445 -465 461
rect -625 411 -609 445
rect -481 411 -465 445
rect -625 364 -465 411
rect -407 445 -247 461
rect -407 411 -391 445
rect -263 411 -247 445
rect -407 364 -247 411
rect -189 445 -29 461
rect -189 411 -173 445
rect -45 411 -29 445
rect -189 364 -29 411
rect 29 445 189 461
rect 29 411 45 445
rect 173 411 189 445
rect 29 364 189 411
rect 247 445 407 461
rect 247 411 263 445
rect 391 411 407 445
rect 247 364 407 411
rect 465 445 625 461
rect 465 411 481 445
rect 609 411 625 445
rect 465 364 625 411
rect 683 445 843 461
rect 683 411 699 445
rect 827 411 843 445
rect 683 364 843 411
rect 901 445 1061 461
rect 901 411 917 445
rect 1045 411 1061 445
rect 901 364 1061 411
rect 1119 445 1279 461
rect 1119 411 1135 445
rect 1263 411 1279 445
rect 1119 364 1279 411
rect -1279 -462 -1119 -436
rect -1061 -462 -901 -436
rect -843 -462 -683 -436
rect -625 -462 -465 -436
rect -407 -462 -247 -436
rect -189 -462 -29 -436
rect 29 -462 189 -436
rect 247 -462 407 -436
rect 465 -462 625 -436
rect 683 -462 843 -436
rect 901 -462 1061 -436
rect 1119 -462 1279 -436
<< polycont >>
rect -1263 411 -1135 445
rect -1045 411 -917 445
rect -827 411 -699 445
rect -609 411 -481 445
rect -391 411 -263 445
rect -173 411 -45 445
rect 45 411 173 445
rect 263 411 391 445
rect 481 411 609 445
rect 699 411 827 445
rect 917 411 1045 445
rect 1135 411 1263 445
<< locali >>
rect -1459 550 -1363 584
rect 1363 550 1459 584
rect -1459 488 -1425 550
rect 1425 488 1459 550
rect -1279 411 -1263 445
rect -1135 411 -1119 445
rect -1061 411 -1045 445
rect -917 411 -901 445
rect -843 411 -827 445
rect -699 411 -683 445
rect -625 411 -609 445
rect -481 411 -465 445
rect -407 411 -391 445
rect -263 411 -247 445
rect -189 411 -173 445
rect -45 411 -29 445
rect 29 411 45 445
rect 173 411 189 445
rect 247 411 263 445
rect 391 411 407 445
rect 465 411 481 445
rect 609 411 625 445
rect 683 411 699 445
rect 827 411 843 445
rect 901 411 917 445
rect 1045 411 1061 445
rect 1119 411 1135 445
rect 1263 411 1279 445
rect -1325 352 -1291 368
rect -1325 -440 -1291 -424
rect -1107 352 -1073 368
rect -1107 -440 -1073 -424
rect -889 352 -855 368
rect -889 -440 -855 -424
rect -671 352 -637 368
rect -671 -440 -637 -424
rect -453 352 -419 368
rect -453 -440 -419 -424
rect -235 352 -201 368
rect -235 -440 -201 -424
rect -17 352 17 368
rect -17 -440 17 -424
rect 201 352 235 368
rect 201 -440 235 -424
rect 419 352 453 368
rect 419 -440 453 -424
rect 637 352 671 368
rect 637 -440 671 -424
rect 855 352 889 368
rect 855 -440 889 -424
rect 1073 352 1107 368
rect 1073 -440 1107 -424
rect 1291 352 1325 368
rect 1291 -440 1325 -424
rect -1459 -550 -1425 -488
rect 1425 -550 1459 -488
rect -1459 -584 -1363 -550
rect 1363 -584 1459 -550
<< viali >>
rect -1263 411 -1135 445
rect -1045 411 -917 445
rect -827 411 -699 445
rect -609 411 -481 445
rect -391 411 -263 445
rect -173 411 -45 445
rect 45 411 173 445
rect 263 411 391 445
rect 481 411 609 445
rect 699 411 827 445
rect 917 411 1045 445
rect 1135 411 1263 445
rect -1325 -424 -1291 352
rect -1107 -424 -1073 352
rect -889 -424 -855 352
rect -671 -424 -637 352
rect -453 -424 -419 352
rect -235 -424 -201 352
rect -17 -424 17 352
rect 201 -424 235 352
rect 419 -424 453 352
rect 637 -424 671 352
rect 855 -424 889 352
rect 1073 -424 1107 352
rect 1291 -424 1325 352
<< metal1 >>
rect -1275 445 -1123 451
rect -1275 411 -1263 445
rect -1135 411 -1123 445
rect -1275 405 -1123 411
rect -1057 445 -905 451
rect -1057 411 -1045 445
rect -917 411 -905 445
rect -1057 405 -905 411
rect -839 445 -687 451
rect -839 411 -827 445
rect -699 411 -687 445
rect -839 405 -687 411
rect -621 445 -469 451
rect -621 411 -609 445
rect -481 411 -469 445
rect -621 405 -469 411
rect -403 445 -251 451
rect -403 411 -391 445
rect -263 411 -251 445
rect -403 405 -251 411
rect -185 445 -33 451
rect -185 411 -173 445
rect -45 411 -33 445
rect -185 405 -33 411
rect 33 445 185 451
rect 33 411 45 445
rect 173 411 185 445
rect 33 405 185 411
rect 251 445 403 451
rect 251 411 263 445
rect 391 411 403 445
rect 251 405 403 411
rect 469 445 621 451
rect 469 411 481 445
rect 609 411 621 445
rect 469 405 621 411
rect 687 445 839 451
rect 687 411 699 445
rect 827 411 839 445
rect 687 405 839 411
rect 905 445 1057 451
rect 905 411 917 445
rect 1045 411 1057 445
rect 905 405 1057 411
rect 1123 445 1275 451
rect 1123 411 1135 445
rect 1263 411 1275 445
rect 1123 405 1275 411
rect -1331 352 -1285 364
rect -1331 -424 -1325 352
rect -1291 -424 -1285 352
rect -1331 -436 -1285 -424
rect -1113 352 -1067 364
rect -1113 -424 -1107 352
rect -1073 -424 -1067 352
rect -1113 -436 -1067 -424
rect -895 352 -849 364
rect -895 -424 -889 352
rect -855 -424 -849 352
rect -895 -436 -849 -424
rect -677 352 -631 364
rect -677 -424 -671 352
rect -637 -424 -631 352
rect -677 -436 -631 -424
rect -459 352 -413 364
rect -459 -424 -453 352
rect -419 -424 -413 352
rect -459 -436 -413 -424
rect -241 352 -195 364
rect -241 -424 -235 352
rect -201 -424 -195 352
rect -241 -436 -195 -424
rect -23 352 23 364
rect -23 -424 -17 352
rect 17 -424 23 352
rect -23 -436 23 -424
rect 195 352 241 364
rect 195 -424 201 352
rect 235 -424 241 352
rect 195 -436 241 -424
rect 413 352 459 364
rect 413 -424 419 352
rect 453 -424 459 352
rect 413 -436 459 -424
rect 631 352 677 364
rect 631 -424 637 352
rect 671 -424 677 352
rect 631 -436 677 -424
rect 849 352 895 364
rect 849 -424 855 352
rect 889 -424 895 352
rect 849 -436 895 -424
rect 1067 352 1113 364
rect 1067 -424 1073 352
rect 1107 -424 1113 352
rect 1067 -436 1113 -424
rect 1285 352 1331 364
rect 1285 -424 1291 352
rect 1325 -424 1331 352
rect 1285 -436 1331 -424
<< properties >>
string FIXED_BBOX -1442 -567 1442 567
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 4 l 0.8 m 1 nf 12 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
