magic
tech sky130a
timestamp 1739287221
<< checkpaint >>
rect -47 -88 757 204
<< l65d20 >>
rect 0 0 710 150
<< l66d44 >>
rect 7 13 24 30
rect 687 13 704 30
rect 7 49 24 66
rect 687 49 704 66
rect 7 85 24 102
rect 687 85 704 102
rect 7 121 24 138
rect 687 121 704 138
rect 347 13 364 30
rect 347 49 364 66
rect 347 85 364 102
rect 347 121 364 138
rect 46 -45 63 -28
rect 396 -45 413 -28
rect 82 -45 99 -28
rect 432 -45 449 -28
rect 118 -45 135 -28
rect 468 -45 485 -28
rect 154 -45 171 -28
rect 504 -45 521 -28
rect 190 -45 207 -28
rect 540 -45 557 -28
rect 226 -45 243 -28
rect 576 -45 593 -28
rect 262 -45 279 -28
rect 612 -45 629 -28
rect 298 -45 315 -28
rect 648 -45 665 -28
<< l67d20 >>
rect 7 5 24 146
rect 687 5 704 146
rect 347 5 364 146
rect 38 -45 323 -28
rect 388 -45 673 -28
<< l67d44 >>
rect 7 13 24 30
rect 687 13 704 30
rect 7 49 24 66
rect 687 49 704 66
rect 7 85 24 102
rect 687 85 704 102
rect 7 121 24 138
rect 687 121 704 138
rect 347 13 364 30
rect 347 49 364 66
rect 347 85 364 102
rect 347 121 364 138
rect 46 -45 63 -28
rect 396 -45 413 -28
rect 82 -45 99 -28
rect 432 -45 449 -28
rect 118 -45 135 -28
rect 468 -45 485 -28
rect 154 -45 171 -28
rect 504 -45 521 -28
rect 190 -45 207 -28
rect 540 -45 557 -28
rect 226 -45 243 -28
rect 576 -45 593 -28
rect 262 -45 279 -28
rect 612 -45 629 -28
rect 298 -45 315 -28
rect 648 -45 665 -28
<< l68d20 >>
rect 4 7 27 144
rect 684 7 707 144
rect 344 7 367 144
rect 40 -48 321 -25
rect 390 -48 671 -25
<< l66d20 >>
rect 30 -53 330 -20
rect 380 -53 680 -20
rect 30 -20 330 170
rect 380 -20 680 170
<< l95d20 >>
rect 29 -54 331 -19
rect 379 -54 681 -19
<< l94d20 >>
rect -13 -13 723 163
<< l64d20 >>
rect -47 -88 757 204
<< l75d20 >>
rect -47 -88 757 204
<< end >>
