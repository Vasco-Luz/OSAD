magic
tech sky130A
magscale 1 2
timestamp 1693700175
<< error_p >>
rect -1228 841 -1170 847
rect -1010 841 -952 847
rect -792 841 -734 847
rect -574 841 -516 847
rect -356 841 -298 847
rect -138 841 -80 847
rect 80 841 138 847
rect 298 841 356 847
rect 516 841 574 847
rect 734 841 792 847
rect 952 841 1010 847
rect 1170 841 1228 847
rect -1228 807 -1216 841
rect -1010 807 -998 841
rect -792 807 -780 841
rect -574 807 -562 841
rect -356 807 -344 841
rect -138 807 -126 841
rect 80 807 92 841
rect 298 807 310 841
rect 516 807 528 841
rect 734 807 746 841
rect 952 807 964 841
rect 1170 807 1182 841
rect -1228 801 -1170 807
rect -1010 801 -952 807
rect -792 801 -734 807
rect -574 801 -516 807
rect -356 801 -298 807
rect -138 801 -80 807
rect 80 801 138 807
rect 298 801 356 807
rect 516 801 574 807
rect 734 801 792 807
rect 952 801 1010 807
rect 1170 801 1228 807
<< pwell >>
rect -1507 -1027 1507 1027
<< mvnmos >>
rect -1279 -831 -1119 769
rect -1061 -831 -901 769
rect -843 -831 -683 769
rect -625 -831 -465 769
rect -407 -831 -247 769
rect -189 -831 -29 769
rect 29 -831 189 769
rect 247 -831 407 769
rect 465 -831 625 769
rect 683 -831 843 769
rect 901 -831 1061 769
rect 1119 -831 1279 769
<< mvndiff >>
rect -1337 757 -1279 769
rect -1337 -819 -1325 757
rect -1291 -819 -1279 757
rect -1337 -831 -1279 -819
rect -1119 757 -1061 769
rect -1119 -819 -1107 757
rect -1073 -819 -1061 757
rect -1119 -831 -1061 -819
rect -901 757 -843 769
rect -901 -819 -889 757
rect -855 -819 -843 757
rect -901 -831 -843 -819
rect -683 757 -625 769
rect -683 -819 -671 757
rect -637 -819 -625 757
rect -683 -831 -625 -819
rect -465 757 -407 769
rect -465 -819 -453 757
rect -419 -819 -407 757
rect -465 -831 -407 -819
rect -247 757 -189 769
rect -247 -819 -235 757
rect -201 -819 -189 757
rect -247 -831 -189 -819
rect -29 757 29 769
rect -29 -819 -17 757
rect 17 -819 29 757
rect -29 -831 29 -819
rect 189 757 247 769
rect 189 -819 201 757
rect 235 -819 247 757
rect 189 -831 247 -819
rect 407 757 465 769
rect 407 -819 419 757
rect 453 -819 465 757
rect 407 -831 465 -819
rect 625 757 683 769
rect 625 -819 637 757
rect 671 -819 683 757
rect 625 -831 683 -819
rect 843 757 901 769
rect 843 -819 855 757
rect 889 -819 901 757
rect 843 -831 901 -819
rect 1061 757 1119 769
rect 1061 -819 1073 757
rect 1107 -819 1119 757
rect 1061 -831 1119 -819
rect 1279 757 1337 769
rect 1279 -819 1291 757
rect 1325 -819 1337 757
rect 1279 -831 1337 -819
<< mvndiffc >>
rect -1325 -819 -1291 757
rect -1107 -819 -1073 757
rect -889 -819 -855 757
rect -671 -819 -637 757
rect -453 -819 -419 757
rect -235 -819 -201 757
rect -17 -819 17 757
rect 201 -819 235 757
rect 419 -819 453 757
rect 637 -819 671 757
rect 855 -819 889 757
rect 1073 -819 1107 757
rect 1291 -819 1325 757
<< mvpsubdiff >>
rect -1471 979 1471 991
rect -1471 945 -1363 979
rect 1363 945 1471 979
rect -1471 933 1471 945
rect -1471 883 -1413 933
rect -1471 -883 -1459 883
rect -1425 -883 -1413 883
rect 1413 883 1471 933
rect -1471 -933 -1413 -883
rect 1413 -883 1425 883
rect 1459 -883 1471 883
rect 1413 -933 1471 -883
rect -1471 -945 1471 -933
rect -1471 -979 -1363 -945
rect 1363 -979 1471 -945
rect -1471 -991 1471 -979
<< mvpsubdiffcont >>
rect -1363 945 1363 979
rect -1459 -883 -1425 883
rect 1425 -883 1459 883
rect -1363 -979 1363 -945
<< poly >>
rect -1232 841 -1166 857
rect -1232 824 -1216 841
rect -1279 807 -1216 824
rect -1182 824 -1166 841
rect -1014 841 -948 857
rect -1014 824 -998 841
rect -1182 807 -1119 824
rect -1279 769 -1119 807
rect -1061 807 -998 824
rect -964 824 -948 841
rect -796 841 -730 857
rect -796 824 -780 841
rect -964 807 -901 824
rect -1061 769 -901 807
rect -843 807 -780 824
rect -746 824 -730 841
rect -578 841 -512 857
rect -578 824 -562 841
rect -746 807 -683 824
rect -843 769 -683 807
rect -625 807 -562 824
rect -528 824 -512 841
rect -360 841 -294 857
rect -360 824 -344 841
rect -528 807 -465 824
rect -625 769 -465 807
rect -407 807 -344 824
rect -310 824 -294 841
rect -142 841 -76 857
rect -142 824 -126 841
rect -310 807 -247 824
rect -407 769 -247 807
rect -189 807 -126 824
rect -92 824 -76 841
rect 76 841 142 857
rect 76 824 92 841
rect -92 807 -29 824
rect -189 769 -29 807
rect 29 807 92 824
rect 126 824 142 841
rect 294 841 360 857
rect 294 824 310 841
rect 126 807 189 824
rect 29 769 189 807
rect 247 807 310 824
rect 344 824 360 841
rect 512 841 578 857
rect 512 824 528 841
rect 344 807 407 824
rect 247 769 407 807
rect 465 807 528 824
rect 562 824 578 841
rect 730 841 796 857
rect 730 824 746 841
rect 562 807 625 824
rect 465 769 625 807
rect 683 807 746 824
rect 780 824 796 841
rect 948 841 1014 857
rect 948 824 964 841
rect 780 807 843 824
rect 683 769 843 807
rect 901 807 964 824
rect 998 824 1014 841
rect 1166 841 1232 857
rect 1166 824 1182 841
rect 998 807 1061 824
rect 901 769 1061 807
rect 1119 807 1182 824
rect 1216 824 1232 841
rect 1216 807 1279 824
rect 1119 769 1279 807
rect -1279 -857 -1119 -831
rect -1061 -857 -901 -831
rect -843 -857 -683 -831
rect -625 -857 -465 -831
rect -407 -857 -247 -831
rect -189 -857 -29 -831
rect 29 -857 189 -831
rect 247 -857 407 -831
rect 465 -857 625 -831
rect 683 -857 843 -831
rect 901 -857 1061 -831
rect 1119 -857 1279 -831
<< polycont >>
rect -1216 807 -1182 841
rect -998 807 -964 841
rect -780 807 -746 841
rect -562 807 -528 841
rect -344 807 -310 841
rect -126 807 -92 841
rect 92 807 126 841
rect 310 807 344 841
rect 528 807 562 841
rect 746 807 780 841
rect 964 807 998 841
rect 1182 807 1216 841
<< locali >>
rect -1459 945 -1363 979
rect 1363 945 1459 979
rect -1459 883 -1425 945
rect 1425 883 1459 945
rect -1232 807 -1216 841
rect -1182 807 -1166 841
rect -1014 807 -998 841
rect -964 807 -948 841
rect -796 807 -780 841
rect -746 807 -730 841
rect -578 807 -562 841
rect -528 807 -512 841
rect -360 807 -344 841
rect -310 807 -294 841
rect -142 807 -126 841
rect -92 807 -76 841
rect 76 807 92 841
rect 126 807 142 841
rect 294 807 310 841
rect 344 807 360 841
rect 512 807 528 841
rect 562 807 578 841
rect 730 807 746 841
rect 780 807 796 841
rect 948 807 964 841
rect 998 807 1014 841
rect 1166 807 1182 841
rect 1216 807 1232 841
rect -1325 757 -1291 773
rect -1325 -835 -1291 -819
rect -1107 757 -1073 773
rect -1107 -835 -1073 -819
rect -889 757 -855 773
rect -889 -835 -855 -819
rect -671 757 -637 773
rect -671 -835 -637 -819
rect -453 757 -419 773
rect -453 -835 -419 -819
rect -235 757 -201 773
rect -235 -835 -201 -819
rect -17 757 17 773
rect -17 -835 17 -819
rect 201 757 235 773
rect 201 -835 235 -819
rect 419 757 453 773
rect 419 -835 453 -819
rect 637 757 671 773
rect 637 -835 671 -819
rect 855 757 889 773
rect 855 -835 889 -819
rect 1073 757 1107 773
rect 1073 -835 1107 -819
rect 1291 757 1325 773
rect 1291 -835 1325 -819
rect -1459 -945 -1425 -883
rect 1425 -945 1459 -883
rect -1459 -979 -1363 -945
rect 1363 -979 1459 -945
<< viali >>
rect -1216 807 -1182 841
rect -998 807 -964 841
rect -780 807 -746 841
rect -562 807 -528 841
rect -344 807 -310 841
rect -126 807 -92 841
rect 92 807 126 841
rect 310 807 344 841
rect 528 807 562 841
rect 746 807 780 841
rect 964 807 998 841
rect 1182 807 1216 841
rect -1325 -819 -1291 757
rect -1107 -819 -1073 757
rect -889 -819 -855 757
rect -671 -819 -637 757
rect -453 -819 -419 757
rect -235 -819 -201 757
rect -17 -819 17 757
rect 201 -819 235 757
rect 419 -819 453 757
rect 637 -819 671 757
rect 855 -819 889 757
rect 1073 -819 1107 757
rect 1291 -819 1325 757
<< metal1 >>
rect -1228 841 -1170 847
rect -1228 807 -1216 841
rect -1182 807 -1170 841
rect -1228 801 -1170 807
rect -1010 841 -952 847
rect -1010 807 -998 841
rect -964 807 -952 841
rect -1010 801 -952 807
rect -792 841 -734 847
rect -792 807 -780 841
rect -746 807 -734 841
rect -792 801 -734 807
rect -574 841 -516 847
rect -574 807 -562 841
rect -528 807 -516 841
rect -574 801 -516 807
rect -356 841 -298 847
rect -356 807 -344 841
rect -310 807 -298 841
rect -356 801 -298 807
rect -138 841 -80 847
rect -138 807 -126 841
rect -92 807 -80 841
rect -138 801 -80 807
rect 80 841 138 847
rect 80 807 92 841
rect 126 807 138 841
rect 80 801 138 807
rect 298 841 356 847
rect 298 807 310 841
rect 344 807 356 841
rect 298 801 356 807
rect 516 841 574 847
rect 516 807 528 841
rect 562 807 574 841
rect 516 801 574 807
rect 734 841 792 847
rect 734 807 746 841
rect 780 807 792 841
rect 734 801 792 807
rect 952 841 1010 847
rect 952 807 964 841
rect 998 807 1010 841
rect 952 801 1010 807
rect 1170 841 1228 847
rect 1170 807 1182 841
rect 1216 807 1228 841
rect 1170 801 1228 807
rect -1331 757 -1285 769
rect -1331 -819 -1325 757
rect -1291 -819 -1285 757
rect -1331 -831 -1285 -819
rect -1113 757 -1067 769
rect -1113 -819 -1107 757
rect -1073 -819 -1067 757
rect -1113 -831 -1067 -819
rect -895 757 -849 769
rect -895 -819 -889 757
rect -855 -819 -849 757
rect -895 -831 -849 -819
rect -677 757 -631 769
rect -677 -819 -671 757
rect -637 -819 -631 757
rect -677 -831 -631 -819
rect -459 757 -413 769
rect -459 -819 -453 757
rect -419 -819 -413 757
rect -459 -831 -413 -819
rect -241 757 -195 769
rect -241 -819 -235 757
rect -201 -819 -195 757
rect -241 -831 -195 -819
rect -23 757 23 769
rect -23 -819 -17 757
rect 17 -819 23 757
rect -23 -831 23 -819
rect 195 757 241 769
rect 195 -819 201 757
rect 235 -819 241 757
rect 195 -831 241 -819
rect 413 757 459 769
rect 413 -819 419 757
rect 453 -819 459 757
rect 413 -831 459 -819
rect 631 757 677 769
rect 631 -819 637 757
rect 671 -819 677 757
rect 631 -831 677 -819
rect 849 757 895 769
rect 849 -819 855 757
rect 889 -819 895 757
rect 849 -831 895 -819
rect 1067 757 1113 769
rect 1067 -819 1073 757
rect 1107 -819 1113 757
rect 1067 -831 1113 -819
rect 1285 757 1331 769
rect 1285 -819 1291 757
rect 1325 -819 1331 757
rect 1285 -831 1331 -819
<< properties >>
string FIXED_BBOX -1442 -962 1442 962
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 8 l 0.8 m 1 nf 12 diffcov 100 polycov 20 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 0.5 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
