** sch_path: /home/vasco/Desktop/sky130A_tests/automatization_analog_design/mos_dc_characteristic/mos.sch
**.subckt mos
V1 net1 GND VD
V2 net2 GND VG
Vmeas net1 net3 0
.save i(vmeas)
XM13 GND net2 net3 GND sky130_fd_pr__pfet_20v0 L=1 W=30 m=1
**** begin user architecture code

**************************************************************
**************************************************************
**************************************************************
**************************************************************
**************************************************************
*LIBs*********************************************************
**************************************************************
**************************************************************
**************************************************************
**************************************************************
**************************************************************
*.lib /home/vasco/PDK/sky130B/libs.tech/ngspice/sky130.lib.spice tt
* chose the corners in the corner file
* tt_mm for mismatch
* ss ff sf fs standart corners
* ll hh lh hl capacitor and resistors corners
* mc for total process variation including corners
**************************************************************
**************************************************************
**************************************************************
**************************************************************
**************************************************************
*Corners/montecarlo options***********************************
**************************************************************
**************************************************************
**************************************************************
**************************************************************
**************************************************************
.TEMP 27
**************************************************************
**************************************************************
**************************************************************
**************************************************************
*SIMULATION and Plots*****************************************
**************************************************************
**************************************************************
**************************************************************
**************************************************************
.control
save all
.endc


.param mc_mm_switch=0
.param mc_pr_switch=0
.include /home/vasco/PDK/sky130B/libs.tech/ngspice/corners/tt.spice
.include /home/vasco/PDK/sky130B/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/vasco/PDK/sky130B/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/vasco/PDK/sky130B/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends
.GLOBAL GND
.end
