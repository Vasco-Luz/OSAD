* Extracted by KLayout with SKY130 LVS runset on : 26/02/2025 00:41

.SUBCKT Pmos_current_mirror
X$1 \$1 vias_gen$2
X$2 \$1 vias_gen
X$3 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1
+ \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1
+ \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1
+ \$1 \$1 \$1 \$1 \$1 \$1 \$1 pfet
X$4 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1
+ \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1
+ \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1 \$1
+ \$1 \$1 \$1 \$1 \$1 \$1 \$1 pfet
X$5 \$1 vias_gen
X$6 \$1 vias_gen
X$7 \$1 vias_gen
X$8 \$1 vias_gen$2
X$9 \$1 vias_gen$2
X$10 \$1 vias_gen$2
X$11 \$1 vias_gen$2
X$12 \$1 vias_gen$2
X$13 \$1 vias_gen$2
X$14 \$1 vias_gen$2
X$15 \$1 vias_gen$2
X$16 \$1 vias_gen$2
X$17 \$1 vias_gen$2
X$18 \$1 vias_gen$2
X$19 \$1 guard_ring_gen$1
.ENDS Pmos_current_mirror

.SUBCKT guard_ring_gen$1 \$1
.ENDS guard_ring_gen$1

.SUBCKT vias_gen$2 \$1
.ENDS vias_gen$2

.SUBCKT pfet \$1 \$2 \$3 \$4 \$5 \$6 \$7 \$8 \$9 \$10 \$11 \$12 \$13 \$14 \$15
+ \$16 \$17 \$18 \$19 \$20 \$21 \$22 \$23 \$24 \$25 \$26 \$27 \$28 \$29 \$30
+ \$31 \$32 \$33 \$34 \$35 \$36 \$37 \$38 \$39 \$40 \$41 \$42 \$43 \$44 \$45
+ \$46 \$47 \$48 \$49 \$50 \$51 \$52 \$53 \$54 \$55 \$56 \$57 \$58 \$59 \$60
+ \$61 \$62 \$63 \$64
M$1 \$32 \$1 \$33 \$64 sky130_fd_pr__pfet_g5v0d10v5 L=2.2 W=1 AS=0.3 AD=0.25
+ PS=2.6 PD=1.5
M$2 \$33 \$2 \$34 \$64 sky130_fd_pr__pfet_g5v0d10v5 L=2.2 W=1 AS=0.25 AD=0.25
+ PS=1.5 PD=1.5
M$3 \$34 \$3 \$35 \$64 sky130_fd_pr__pfet_g5v0d10v5 L=2.2 W=1 AS=0.25 AD=0.25
+ PS=1.5 PD=1.5
M$4 \$35 \$4 \$36 \$64 sky130_fd_pr__pfet_g5v0d10v5 L=2.2 W=1 AS=0.25 AD=0.25
+ PS=1.5 PD=1.5
M$5 \$36 \$5 \$37 \$64 sky130_fd_pr__pfet_g5v0d10v5 L=2.2 W=1 AS=0.25 AD=0.25
+ PS=1.5 PD=1.5
M$6 \$37 \$6 \$38 \$64 sky130_fd_pr__pfet_g5v0d10v5 L=2.2 W=1 AS=0.25 AD=0.25
+ PS=1.5 PD=1.5
M$7 \$38 \$7 \$39 \$64 sky130_fd_pr__pfet_g5v0d10v5 L=2.2 W=1 AS=0.25 AD=0.25
+ PS=1.5 PD=1.5
M$8 \$39 \$8 \$40 \$64 sky130_fd_pr__pfet_g5v0d10v5 L=2.2 W=1 AS=0.25 AD=0.25
+ PS=1.5 PD=1.5
M$9 \$40 \$9 \$41 \$64 sky130_fd_pr__pfet_g5v0d10v5 L=2.2 W=1 AS=0.25 AD=0.25
+ PS=1.5 PD=1.5
M$10 \$41 \$10 \$42 \$64 sky130_fd_pr__pfet_g5v0d10v5 L=2.2 W=1 AS=0.25 AD=0.25
+ PS=1.5 PD=1.5
M$11 \$42 \$11 \$43 \$64 sky130_fd_pr__pfet_g5v0d10v5 L=2.2 W=1 AS=0.25 AD=0.25
+ PS=1.5 PD=1.5
M$12 \$43 \$12 \$44 \$64 sky130_fd_pr__pfet_g5v0d10v5 L=2.2 W=1 AS=0.25 AD=0.25
+ PS=1.5 PD=1.5
M$13 \$44 \$13 \$45 \$64 sky130_fd_pr__pfet_g5v0d10v5 L=2.2 W=1 AS=0.25 AD=0.25
+ PS=1.5 PD=1.5
M$14 \$45 \$14 \$46 \$64 sky130_fd_pr__pfet_g5v0d10v5 L=2.2 W=1 AS=0.25 AD=0.25
+ PS=1.5 PD=1.5
M$15 \$46 \$15 \$47 \$64 sky130_fd_pr__pfet_g5v0d10v5 L=2.2 W=1 AS=0.25 AD=0.25
+ PS=1.5 PD=1.5
M$16 \$47 \$16 \$48 \$64 sky130_fd_pr__pfet_g5v0d10v5 L=2.2 W=1 AS=0.25 AD=0.25
+ PS=1.5 PD=1.5
M$17 \$48 \$17 \$49 \$64 sky130_fd_pr__pfet_g5v0d10v5 L=2.2 W=1 AS=0.25 AD=0.25
+ PS=1.5 PD=1.5
M$18 \$49 \$18 \$50 \$64 sky130_fd_pr__pfet_g5v0d10v5 L=2.2 W=1 AS=0.25 AD=0.25
+ PS=1.5 PD=1.5
M$19 \$50 \$19 \$51 \$64 sky130_fd_pr__pfet_g5v0d10v5 L=2.2 W=1 AS=0.25 AD=0.25
+ PS=1.5 PD=1.5
M$20 \$51 \$20 \$52 \$64 sky130_fd_pr__pfet_g5v0d10v5 L=2.2 W=1 AS=0.25 AD=0.25
+ PS=1.5 PD=1.5
M$21 \$52 \$21 \$53 \$64 sky130_fd_pr__pfet_g5v0d10v5 L=2.2 W=1 AS=0.25 AD=0.25
+ PS=1.5 PD=1.5
M$22 \$53 \$22 \$54 \$64 sky130_fd_pr__pfet_g5v0d10v5 L=2.2 W=1 AS=0.25 AD=0.25
+ PS=1.5 PD=1.5
M$23 \$54 \$23 \$55 \$64 sky130_fd_pr__pfet_g5v0d10v5 L=2.2 W=1 AS=0.25 AD=0.25
+ PS=1.5 PD=1.5
M$24 \$55 \$24 \$56 \$64 sky130_fd_pr__pfet_g5v0d10v5 L=2.2 W=1 AS=0.25 AD=0.25
+ PS=1.5 PD=1.5
M$25 \$56 \$25 \$57 \$64 sky130_fd_pr__pfet_g5v0d10v5 L=2.2 W=1 AS=0.25 AD=0.25
+ PS=1.5 PD=1.5
M$26 \$57 \$26 \$58 \$64 sky130_fd_pr__pfet_g5v0d10v5 L=2.2 W=1 AS=0.25 AD=0.25
+ PS=1.5 PD=1.5
M$27 \$58 \$27 \$59 \$64 sky130_fd_pr__pfet_g5v0d10v5 L=2.2 W=1 AS=0.25 AD=0.25
+ PS=1.5 PD=1.5
M$28 \$59 \$28 \$60 \$64 sky130_fd_pr__pfet_g5v0d10v5 L=2.2 W=1 AS=0.25 AD=0.25
+ PS=1.5 PD=1.5
M$29 \$60 \$29 \$61 \$64 sky130_fd_pr__pfet_g5v0d10v5 L=2.2 W=1 AS=0.25 AD=0.25
+ PS=1.5 PD=1.5
M$30 \$61 \$30 \$62 \$64 sky130_fd_pr__pfet_g5v0d10v5 L=2.2 W=1 AS=0.25 AD=0.25
+ PS=1.5 PD=1.5
M$31 \$62 \$31 \$63 \$64 sky130_fd_pr__pfet_g5v0d10v5 L=2.2 W=1 AS=0.25 AD=0.3
+ PS=1.5 PD=2.6
.ENDS pfet

.SUBCKT vias_gen \$1
.ENDS vias_gen
