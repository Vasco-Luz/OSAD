** sch_path: /home/vasco/Desktop/sky130A_tests/automatization_analog_design/mos_dc_characteristic/mos.sch
**.subckt mos
Vmeas net1 net3 0
XM1 net1 net2 net3 net4 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
**** begin user architecture code

**************************************************************
**************************************************************
**************************************************************
**************************************************************
**************************************************************
*LIBs*********************************************************
**************************************************************
**************************************************************
**************************************************************
**************************************************************
**************************************************************
*.lib /home/vasco/PDK/sky130B/libs.tech/ngspice/sky130.lib.spice tt
* chose the corners in the corner file
* tt_mm for mismatch
* ss ff sf fs standart corners
* ll hh lh hl capacitor and resistors corners
* mc for total process variation including corners
**************************************************************
**************************************************************
**************************************************************
**************************************************************
**************************************************************
*Corners/montecarlo options***********************************
**************************************************************
**************************************************************
**************************************************************
**************************************************************
**************************************************************
.TEMP 27
**************************************************************
**************************************************************
**************************************************************
**************************************************************
*SIMULATION and Plots*****************************************
**************************************************************
**************************************************************
**************************************************************
**************************************************************
.control
save all
.endc


.param mc_mm_switch=0
.param mc_pr_switch=0
.include /home/vasco/PDK/sky130B/libs.tech/ngspice/corners/tt.spice
.include /home/vasco/PDK/sky130B/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/vasco/PDK/sky130B/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/vasco/PDK/sky130B/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends
.end
