** sch_path: /foss/designs/OSAD/Learning/single_ended_amplifiers/two_stage_OTA_testing_scripts/amplifier_design/OTA_mc_ac_tb.sch
**.subckt OTA_mc_ac_tb
V1 VDD GND VDD
V2 VSS GND VSS
Vmeas VDD net2 0
.save i(vmeas)
x1 net2 VSS Va VIN+ VOUT UUT_VA_sky
C1 VOUT VSS CL m=1
V5 net1 GND VCM
V3 VIN+ net1 ac 0.5
V4 net3 VSS ac -0.5
E1 Va net3 net4 VSS 1
R1 VOUT net4 1k ac=1000000000000G m=1
C2 net4 VSS 3p m=1
x2 VDD net17 net7 net6 VOUT_CM UUT_VA_sky
C3 VOUT_CM VSS CL m=1
V7 net5 GND ac 1
E2 net7 net5 net8 VSS 1
R2 VOUT_CM net8 1k ac=1000000000000G m=1
C4 net8 VSS 3p m=1
x3 VDD net12 net10 net9 VOUT_A- UUT_VA_sky
C5 VOUT_A- VSS CL m=1
E3 net10 GND net11 VSS 1
R3 VOUT_A- net11 1k ac=1000000000000G m=1
C6 net11 VSS 3p m=1
V9 net12 VSS ac 1
x4 net13 VSS net15 net14 VOUT_A+ UUT_VA_sky
C7 VOUT_A+ VSS CL m=1
E4 net15 GND net16 VSS 1
R4 VOUT_A+ net16 1k ac=1000000000000G m=1
C8 net16 VSS 3p m=1
V11 net13 VDD ac 1
V8 net9 GND VCM
V12 net14 GND VCM
V6 net6 net5 VCM
**** begin user architecture code
.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice mc

.Temp 27
.param VDD = 5
.param VSS = 0
.param CL = 3p
.param VCM = 2.5
.param mc_mm_switch = 1


.control

	save all
	ac dec 100 1 10G
	plot db(v(VOUT))
	plot db(v(VOUT_CM))
	plot db(v(VOUT_A-))
	plot db(v(VOUT_A+))
	wrdata mc_ac.csv db(v(VOUT)) phase(v(VOUT)) db(v(VOUT_CM)) db(v(VOUT_A-)) db(v(VOUT_A+))
	noise v(VOUT,VSS) V3 dec 10 1 10G
	setplot noise1

	plot onoise_spectrum inoise_spectrum

.endc


**** end user architecture code
**.ends

* expanding   symbol:  Sky130A/UUT_sky/UUT_VA_sky.sym # of pins=5
** sym_path: /foss/designs/OSAD/LIB/Sky130A/UUT_sky/UUT_VA_sky.sym
** sch_path: /foss/designs/OSAD/LIB/Sky130A/UUT_sky/UUT_VA_sky.sch
.subckt UUT_VA_sky VDD VSS VIN- VIN+ VOUT
*.iopin VDD
*.iopin VSS
*.iopin VIN-
*.iopin VIN+
*.iopin VOUT
x1 VDD VSS VIN+ VIN- VOUT VA001_sky130_1_8V
.ends


* expanding   symbol:  Sky130A/single ended amplifiers/VA001_sky130_1_8V.sym # of pins=5
** sym_path: /foss/designs/OSAD/LIB/Sky130A/single ended amplifiers/VA001_sky130_1_8V.sym
** sch_path: /foss/designs/OSAD/LIB/Sky130A/single ended amplifiers/VA001_sky130_1_8V.sch
.subckt VA001_sky130_1_8V VDD VSS Vin+ Vin- VOUT
*.iopin VDD
*.iopin VSS
*.iopin Vin+
*.iopin Vin-
*.iopin VOUT
XR6 VSS net3 VSS sky130_fd_pr__res_high_po_0p35 L=16 mult=1 m=1
XM1 net1 net2 net3 VSS sky130_fd_pr__nfet_01v8 L=4 W='1 * 8 ' nf=8 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=2
+ m=2
XM2 net2 net2 VSS VSS sky130_fd_pr__nfet_01v8 L=4 W='1 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=2
+ m=2
XM5 VB1 VB1 VDD VDD sky130_fd_pr__pfet_01v8 L=2 W='1 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=2
+ m=2
XM6 VB2 VB1 VDD VDD sky130_fd_pr__pfet_01v8 L=2 W='1 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=2
+ m=2
XM7 net4 VB1 VDD VDD sky130_fd_pr__pfet_01v8 L=2 W='1 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=8
+ m=8
XM10 net5 net5 VSS VSS sky130_fd_pr__nfet_01v8 L=2 W='2.3 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=2
+ m=2
XM11 net6 net5 VSS VSS sky130_fd_pr__nfet_01v8 L=2 W='2.3 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=2
+ m=2
XM12 VOUT VB1 VDD VDD sky130_fd_pr__pfet_01v8 L=2 W='1 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=16
+ m=16
XM14 net7 VB2 net6 VSS sky130_fd_pr__nfet_01v8 L=1.9 W='2 * 1 ' nf=1 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=2
+ m=2
XC1 VOUT net7 sky130_fd_pr__cap_mim_m3_1 W=7.6 L=7.6 MF=4 m=4
XM8 net5 Vin- net4 net4 sky130_fd_pr__pfet_01v8_lvt L=0.8 W='2 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=4
+ m=4
XM9 net6 Vin+ net4 net4 sky130_fd_pr__pfet_01v8_lvt L=0.8 W='2 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=4
+ m=4
XM33 VOUT net6 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.5 W='1.5 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=2
+ m=2
XM3 VB2 VB2 net2 VSS sky130_fd_pr__nfet_01v8_lvt L=2 W='1 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=2
+ m=2
XM4 VB1 VB2 net1 VSS sky130_fd_pr__nfet_01v8_lvt L=2 W='1 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=2
+ m=2
.ends

.GLOBAL GND
.end
