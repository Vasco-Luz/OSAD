magic
tech sky130A
magscale 1 2
timestamp 1740482431
<< mvnmos >>
rect -50 -73 50 11
<< mvndiff >>
rect -108 -1 -50 11
rect -108 -61 -96 -1
rect -62 -61 -50 -1
rect -108 -73 -50 -61
rect 50 -1 108 11
rect 50 -61 62 -1
rect 96 -61 108 -1
rect 50 -73 108 -61
<< mvndiffc >>
rect -96 -61 -62 -1
rect 62 -61 96 -1
<< poly >>
rect -43 83 43 99
rect -43 66 -27 83
rect -50 49 -27 66
rect 27 66 43 83
rect 27 49 50 66
rect -50 11 50 49
rect -50 -99 50 -73
<< polycont >>
rect -27 49 27 83
<< locali >>
rect -43 49 -27 83
rect 27 49 43 83
rect -96 -1 -62 15
rect -96 -77 -62 -61
rect 62 -1 96 15
rect 62 -77 96 -61
<< viali >>
rect -27 49 27 83
rect -96 -61 -62 -1
rect 62 -61 96 -1
<< metal1 >>
rect -39 83 39 89
rect -39 49 -27 83
rect 27 49 39 83
rect -39 43 39 49
rect -102 -1 -56 11
rect -102 -61 -96 -1
rect -62 -61 -56 -1
rect -102 -73 -56 -61
rect 56 -1 102 11
rect 56 -61 62 -1
rect 96 -61 102 -1
rect 56 -73 102 -61
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 0.420 l 0.50 m 1 nf 1 diffcov 100 polycov 80 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 80 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
