magic
tech gf180mcuD
magscale 1 10
timestamp 1714262332
<< error_p >>
rect -34 4381 -23 4427
rect 23 4381 34 4392
rect -80 2350 -59 2361
rect 59 2350 80 2361
rect -34 2269 -23 2315
rect -34 2149 -23 2195
rect 23 2149 34 2160
rect -80 118 -59 129
rect 59 118 80 129
rect -34 37 -23 83
rect -34 -83 -23 -37
rect 23 -83 34 -72
rect -80 -2114 -59 -2103
rect 59 -2114 80 -2103
rect -34 -2195 -23 -2149
rect -34 -2315 -23 -2269
rect 23 -2315 34 -2304
rect -80 -4346 -59 -4335
rect 59 -4346 80 -4335
rect -34 -4427 -23 -4381
<< nwell >>
rect -280 -4558 280 4558
<< pmos >>
rect -30 2348 30 4348
rect -30 116 30 2116
rect -30 -2116 30 -116
rect -30 -4348 30 -2348
<< pdiff >>
rect -118 4335 -30 4348
rect -118 2361 -105 4335
rect -59 2361 -30 4335
rect -118 2348 -30 2361
rect 30 4335 118 4348
rect 30 2361 59 4335
rect 105 2361 118 4335
rect 30 2348 118 2361
rect -118 2103 -30 2116
rect -118 129 -105 2103
rect -59 129 -30 2103
rect -118 116 -30 129
rect 30 2103 118 2116
rect 30 129 59 2103
rect 105 129 118 2103
rect 30 116 118 129
rect -118 -129 -30 -116
rect -118 -2103 -105 -129
rect -59 -2103 -30 -129
rect -118 -2116 -30 -2103
rect 30 -129 118 -116
rect 30 -2103 59 -129
rect 105 -2103 118 -129
rect 30 -2116 118 -2103
rect -118 -2361 -30 -2348
rect -118 -4335 -105 -2361
rect -59 -4335 -30 -2361
rect -118 -4348 -30 -4335
rect 30 -2361 118 -2348
rect 30 -4335 59 -2361
rect 105 -4335 118 -2361
rect 30 -4348 118 -4335
<< pdiffc >>
rect -105 2361 -59 4335
rect 59 2361 105 4335
rect -105 129 -59 2103
rect 59 129 105 2103
rect -105 -2103 -59 -129
rect 59 -2103 105 -129
rect -105 -4335 -59 -2361
rect 59 -4335 105 -2361
<< nsubdiff >>
rect -256 4462 256 4534
rect -256 4418 -184 4462
rect -256 -4418 -243 4418
rect -197 -4418 -184 4418
rect 184 4418 256 4462
rect -256 -4462 -184 -4418
rect 184 -4418 197 4418
rect 243 -4418 256 4418
rect 184 -4462 256 -4418
rect -256 -4534 256 -4462
<< nsubdiffcont >>
rect -243 -4418 -197 4418
rect 197 -4418 243 4418
<< polysilicon >>
rect -36 4427 36 4440
rect -36 4381 -23 4427
rect 23 4381 36 4427
rect -36 4368 36 4381
rect -30 4348 30 4368
rect -30 2328 30 2348
rect -36 2315 36 2328
rect -36 2269 -23 2315
rect 23 2269 36 2315
rect -36 2256 36 2269
rect -36 2195 36 2208
rect -36 2149 -23 2195
rect 23 2149 36 2195
rect -36 2136 36 2149
rect -30 2116 30 2136
rect -30 96 30 116
rect -36 83 36 96
rect -36 37 -23 83
rect 23 37 36 83
rect -36 24 36 37
rect -36 -37 36 -24
rect -36 -83 -23 -37
rect 23 -83 36 -37
rect -36 -96 36 -83
rect -30 -116 30 -96
rect -30 -2136 30 -2116
rect -36 -2149 36 -2136
rect -36 -2195 -23 -2149
rect 23 -2195 36 -2149
rect -36 -2208 36 -2195
rect -36 -2269 36 -2256
rect -36 -2315 -23 -2269
rect 23 -2315 36 -2269
rect -36 -2328 36 -2315
rect -30 -2348 30 -2328
rect -30 -4368 30 -4348
rect -36 -4381 36 -4368
rect -36 -4427 -23 -4381
rect 23 -4427 36 -4381
rect -36 -4440 36 -4427
<< polycontact >>
rect -23 4381 23 4427
rect -23 2269 23 2315
rect -23 2149 23 2195
rect -23 37 23 83
rect -23 -83 23 -37
rect -23 -2195 23 -2149
rect -23 -2315 23 -2269
rect -23 -4427 23 -4381
<< metal1 >>
rect -243 4475 243 4521
rect -243 4418 -197 4475
rect -34 4381 -23 4427
rect 23 4381 34 4427
rect 197 4418 243 4475
rect -105 4335 -59 4346
rect -105 2350 -59 2361
rect 59 4335 105 4346
rect 59 2350 105 2361
rect -34 2269 -23 2315
rect 23 2269 34 2315
rect -34 2149 -23 2195
rect 23 2149 34 2195
rect -105 2103 -59 2114
rect -105 118 -59 129
rect 59 2103 105 2114
rect 59 118 105 129
rect -34 37 -23 83
rect 23 37 34 83
rect -34 -83 -23 -37
rect 23 -83 34 -37
rect -105 -129 -59 -118
rect -105 -2114 -59 -2103
rect 59 -129 105 -118
rect 59 -2114 105 -2103
rect -34 -2195 -23 -2149
rect 23 -2195 34 -2149
rect -34 -2315 -23 -2269
rect 23 -2315 34 -2269
rect -105 -2361 -59 -2350
rect -105 -4346 -59 -4335
rect 59 -2361 105 -2350
rect 59 -4346 105 -4335
rect -243 -4475 -197 -4418
rect -34 -4427 -23 -4381
rect 23 -4427 34 -4381
rect 197 -4475 243 -4418
rect -243 -4521 243 -4475
<< properties >>
string FIXED_BBOX -220 -4498 220 4498
string gencell pfet_03v3
string library gf180mcu
string parameters w 10.0 l 0.3 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 1 compatible {pfet_03v3 pfet_06v0}
<< end >>
