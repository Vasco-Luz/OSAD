* NGSPICE file created from TOP.ext - technology: sky130A

.subckt pmos_current_mirror VDD IB IA
X0 IA VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.45 pd=3.6 as=0.45 ps=3.6 w=1.5 l=3
X1 VDD VDD IA VDD sky130_fd_pr__pfet_g5v0d10v5 ad=3.60002 pd=28.805 as=1.80002 ps=14.405 w=1.5 l=3
X2 VDD VDD IA VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1.5 l=3
X3 IA IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1.5 l=3
X4 IA VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1.5 l=3
X5 IA IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1.5 l=3
X6 VDD IA IA VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1.5 l=3
X7 VDD IA IA VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1.5 l=3
X8 VDD IA IB VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.45 pd=3.6 as=0.375 ps=2 w=1.5 l=3
X9 IB IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.375 pd=2 as=0.45 ps=3.6 w=1.5 l=3
X10 VDD IA IB VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=1.5 ps=8 w=1.5 l=3
X11 IB IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1.5 l=3
C0 VDD IA 8.63977f
C1 IA VSUBS 5.0778f
C2 VDD VSUBS 25.41407f
.ends
