magic
tech sky130A
magscale 1 2
timestamp 1740410531
<< nwell >>
rect -273 -1395 2859 1227
<< mvnsubdiff >>
rect -207 1127 -147 1161
rect 2733 1127 2793 1161
rect -207 1101 -173 1127
rect -207 -1295 -173 -1269
rect 2759 1101 2793 1127
rect 2759 -1295 2793 -1269
rect -207 -1329 -147 -1295
rect 2733 -1329 2793 -1295
<< mvnsubdiffcont >>
rect -147 1127 2733 1161
rect -207 -1269 -173 1101
rect 2759 -1269 2793 1101
rect -147 -1329 2733 -1295
<< locali >>
rect -286 1244 2854 1246
rect -286 1238 2968 1244
rect -446 1161 2968 1238
rect -446 1127 -147 1161
rect 2733 1127 2968 1161
rect -446 1116 2968 1127
rect -446 1101 -164 1116
rect -446 -1260 -207 1101
rect -462 -1269 -207 -1260
rect -173 -1260 -164 1101
rect 2740 1101 2968 1116
rect 2740 -1260 2759 1101
rect -173 -1269 2759 -1260
rect 2793 -1260 2968 1101
rect 2793 -1269 2972 -1260
rect -462 -1295 2972 -1269
rect -462 -1329 -147 -1295
rect 2733 -1329 2972 -1295
rect -462 -1418 2972 -1329
<< metal1 >>
rect 3144 1452 3208 1458
rect 3144 1400 3150 1452
rect 3202 1400 3208 1452
rect 3144 1358 3208 1400
rect 3030 1328 3094 1334
rect 3030 1276 3036 1328
rect 3088 1276 3094 1328
rect 3144 1306 3150 1358
rect 3202 1306 3208 1358
rect 3144 1300 3208 1306
rect 3030 1234 3094 1276
rect 3030 1182 3036 1234
rect 3088 1182 3094 1234
rect 3030 1176 3094 1182
rect 3036 -1556 3088 1176
rect 3150 -1358 3202 1300
rect 3144 -1364 3208 -1358
rect 3144 -1416 3150 -1364
rect 3202 -1416 3208 -1364
rect 3144 -1458 3208 -1416
rect 3144 -1510 3150 -1458
rect 3202 -1510 3208 -1458
rect 3144 -1516 3208 -1510
rect 3032 -1562 3096 -1556
rect 3032 -1614 3038 -1562
rect 3090 -1614 3096 -1562
rect 3032 -1656 3096 -1614
rect 3032 -1708 3038 -1656
rect 3090 -1708 3096 -1656
rect 3032 -1714 3096 -1708
<< via1 >>
rect 3150 1400 3202 1452
rect 3036 1276 3088 1328
rect 3150 1306 3202 1358
rect 3036 1182 3088 1234
rect 3150 -1416 3202 -1364
rect 3150 -1510 3202 -1458
rect 3038 -1614 3090 -1562
rect 3038 -1708 3090 -1656
<< metal2 >>
rect 1298 1452 3208 1458
rect 1298 1400 3150 1452
rect 3202 1400 3208 1452
rect 3144 1358 3208 1400
rect 606 1328 3094 1334
rect 606 1280 3036 1328
rect 3030 1276 3036 1280
rect 3088 1276 3094 1328
rect 3144 1306 3150 1358
rect 3202 1306 3208 1358
rect 3144 1300 3208 1306
rect 3030 1234 3094 1276
rect 3030 1182 3036 1234
rect 3088 1182 3094 1234
rect 3030 1176 3094 1182
rect -534 -66 520 -38
rect -588 -146 300 -118
rect 3144 -1364 3208 -1358
rect 3144 -1416 3150 -1364
rect 3202 -1416 3208 -1364
rect 3144 -1458 3208 -1416
rect 3144 -1464 3150 -1458
rect 512 -1510 3150 -1464
rect 3202 -1510 3208 -1458
rect 512 -1516 3208 -1510
rect 3032 -1562 3096 -1556
rect 3032 -1584 3038 -1562
rect 1396 -1614 3038 -1584
rect 3090 -1614 3096 -1562
rect 1396 -1636 3096 -1614
rect 3032 -1656 3096 -1636
rect 3032 -1708 3038 -1656
rect 3090 -1708 3096 -1656
rect 3032 -1714 3096 -1708
use sky130_fd_pr__pfet_g5v0d10v5_AEQKCY  sky130_fd_pr__pfet_g5v0d10v5_AEQKCY_0
timestamp 1740408349
transform 1 0 134 0 -1 -690
box -224 -514 224 640
use sky130_fd_pr__pfet_g5v0d10v5_AEQKCY  sky130_fd_pr__pfet_g5v0d10v5_AEQKCY_1
timestamp 1740408349
transform -1 0 2456 0 -1 -690
box -224 -514 224 640
use sky130_fd_pr__pfet_g5v0d10v5_AEQKCY  sky130_fd_pr__pfet_g5v0d10v5_AEQKCY_2
timestamp 1740408349
transform 1 0 134 0 1 506
box -224 -514 224 640
use sky130_fd_pr__pfet_g5v0d10v5_AEQKCY  sky130_fd_pr__pfet_g5v0d10v5_AEQKCY_3
timestamp 1740408349
transform -1 0 2456 0 1 506
box -224 -514 224 640
use sky130_fd_pr__pfet_g5v0d10v5_PDQKC8  sky130_fd_pr__pfet_g5v0d10v5_PDQKC8_0
timestamp 1740409548
transform -1 0 1295 0 -1 -690
box -645 -596 675 952
use sky130_fd_pr__pfet_g5v0d10v5_PDQKC8  sky130_fd_pr__pfet_g5v0d10v5_PDQKC8_1
timestamp 1740409548
transform 1 0 1295 0 1 506
box -645 -596 675 952
use sky130_fd_pr__pfet_g5v0d10v5_QCQKCQ  sky130_fd_pr__pfet_g5v0d10v5_QCQKCQ_0
timestamp 1740409401
transform -1 0 521 0 -1 -690
box -353 -666 353 832
use sky130_fd_pr__pfet_g5v0d10v5_QCQKCQ  sky130_fd_pr__pfet_g5v0d10v5_QCQKCQ_1
timestamp 1740409401
transform 1 0 2069 0 -1 -690
box -353 -666 353 832
use sky130_fd_pr__pfet_g5v0d10v5_QCQKCQ  sky130_fd_pr__pfet_g5v0d10v5_QCQKCQ_2
timestamp 1740409401
transform 1 0 521 0 1 506
box -353 -666 353 832
use sky130_fd_pr__pfet_g5v0d10v5_QCQKCQ  sky130_fd_pr__pfet_g5v0d10v5_QCQKCQ_3
timestamp 1740409401
transform -1 0 2069 0 1 506
box -353 -666 353 832
<< labels >>
flabel metal2 -574 -136 -548 -126 0 FreeSans 1600 0 0 0 Vin+
port 5 nsew
flabel metal2 -508 -62 -496 -40 0 FreeSans 1600 0 0 0 Vin-
port 7 nsew
flabel locali -386 1066 -306 1188 0 FreeSans 1600 0 0 0 Ibias
port 9 nsew
flabel metal2 720 -1500 750 -1484 0 FreeSans 1600 0 0 0 Ia
port 11 nsew
flabel metal2 1746 -1624 1822 -1594 0 FreeSans 1600 0 0 0 Ib
port 13 nsew
<< end >>
