magic
tech sky130A
magscale 1 2
timestamp 1730492473
<< nwell >>
rect -2802 624 1275 786
<< poly >>
rect -2709 609 -2109 697
rect -2709 569 -2540 609
rect -2270 569 -2109 609
rect -2709 547 -2109 569
rect -2051 602 -1451 697
rect -2051 562 -1882 602
rect -1612 562 -1451 602
rect -2051 540 -1451 562
rect -1393 608 -793 697
rect -1393 568 -1224 608
rect -954 568 -793 608
rect -1393 546 -793 568
rect -735 601 -135 697
rect -735 561 -566 601
rect -296 561 -135 601
rect -735 539 -135 561
rect -77 608 523 697
rect -77 568 92 608
rect 362 568 523 608
rect -77 546 523 568
rect 581 601 1181 697
rect 581 561 750 601
rect 1020 561 1181 601
rect 581 539 1181 561
<< polycont >>
rect -2540 569 -2270 609
rect -1882 562 -1612 602
rect -1224 568 -954 608
rect -566 561 -296 601
rect 92 568 362 608
rect 750 561 1020 601
<< locali >>
rect -2556 609 -2254 625
rect -2556 569 -2540 609
rect -2270 569 -2254 609
rect -2556 551 -2254 569
rect -1898 602 -1596 618
rect -1898 562 -1882 602
rect -1612 562 -1596 602
rect -1898 544 -1596 562
rect -1240 608 -938 624
rect -1240 568 -1224 608
rect -954 568 -938 608
rect -1240 550 -938 568
rect -582 601 -280 617
rect -582 561 -566 601
rect -296 561 -280 601
rect -582 543 -280 561
rect 76 608 378 624
rect 76 568 92 608
rect 362 568 378 608
rect 76 550 378 568
rect 734 601 1036 617
rect 734 561 750 601
rect 1020 561 1036 601
rect 734 543 1036 561
<< viali >>
rect -2540 569 -2270 609
rect -1882 562 -1612 602
rect -1224 568 -954 608
rect -566 561 -296 601
rect 92 568 362 608
rect 750 561 1020 601
<< metal1 >>
rect -2556 619 -2254 639
rect -2556 567 -2540 619
rect -2270 567 -2254 619
rect -2556 551 -2254 567
rect -1898 612 -1596 632
rect -1898 560 -1882 612
rect -1612 560 -1596 612
rect -1898 544 -1596 560
rect -1240 618 -938 638
rect -1240 566 -1224 618
rect -954 566 -938 618
rect -1240 550 -938 566
rect -582 611 -280 631
rect -582 559 -566 611
rect -296 559 -280 611
rect -582 543 -280 559
rect 76 618 378 638
rect 76 566 92 618
rect 362 566 378 618
rect 76 550 378 566
rect 734 611 1036 631
rect 734 559 750 611
rect 1020 559 1036 611
rect 734 543 1036 559
<< via1 >>
rect -2540 609 -2270 619
rect -2540 569 -2270 609
rect -2540 567 -2270 569
rect -1882 602 -1612 612
rect -1882 562 -1612 602
rect -1882 560 -1612 562
rect -1224 608 -954 618
rect -1224 568 -954 608
rect -1224 566 -954 568
rect -566 601 -296 611
rect -566 561 -296 601
rect -566 559 -296 561
rect 92 608 362 618
rect 92 568 362 608
rect 92 566 362 568
rect 750 601 1020 611
rect 750 561 1020 601
rect 750 559 1020 561
<< metal2 >>
rect -2556 625 -2254 629
rect -2556 567 -2540 625
rect -2270 567 -2254 625
rect -1240 624 -938 628
rect -2556 551 -2254 567
rect -1898 618 -1596 622
rect -1898 560 -1882 618
rect -1612 560 -1596 618
rect -1898 544 -1596 560
rect -1240 566 -1224 624
rect -954 566 -938 624
rect 76 624 378 628
rect -1240 550 -938 566
rect -582 617 -280 621
rect -582 559 -566 617
rect -296 559 -280 617
rect -582 543 -280 559
rect 76 566 92 624
rect 362 566 378 624
rect 76 550 378 566
rect 734 617 1036 621
rect 734 559 750 617
rect 1020 559 1036 617
rect 734 543 1036 559
<< via2 >>
rect -2540 619 -2270 625
rect -2540 569 -2270 619
rect -1882 612 -1612 618
rect -1882 562 -1612 612
rect -1224 618 -954 624
rect -1224 568 -954 618
rect -566 611 -296 617
rect -566 561 -296 611
rect 92 618 362 624
rect 92 568 362 618
rect 750 611 1020 617
rect 750 561 1020 611
<< metal3 >>
rect -2556 625 -2254 633
rect -2556 569 -2540 625
rect -2270 569 -2254 625
rect -2556 551 -2254 569
rect -1898 618 -1596 626
rect -1898 562 -1882 618
rect -1612 562 -1596 618
rect -1898 544 -1596 562
rect -1240 624 -938 632
rect -1240 568 -1224 624
rect -954 568 -938 624
rect -1240 550 -938 568
rect -582 617 -280 625
rect -582 561 -566 617
rect -296 561 -280 617
rect -582 543 -280 561
rect 76 624 378 632
rect 76 568 92 624
rect 362 568 378 624
rect 76 550 378 568
rect 734 617 1036 625
rect 734 561 750 617
rect 1020 561 1036 617
rect 734 543 1036 561
use sky130_fd_pr__pfet_01v8_455LYC  sky130_fd_pr__pfet_01v8_455LYC_0 ~/Desktop/OSAD/my_ip/Layouts/VA001_PMOS_1.8_sky130
timestamp 1730491634
transform 1 0 223 0 1 1123
box -394 -462 394 462
use sky130_fd_pr__pfet_01v8_455LYC  sky130_fd_pr__pfet_01v8_455LYC_1
timestamp 1730491634
transform 1 0 -1093 0 1 1123
box -394 -462 394 462
use sky130_fd_pr__pfet_01v8_455LYC  sky130_fd_pr__pfet_01v8_455LYC_2
timestamp 1730491634
transform 1 0 -1751 0 1 1123
box -394 -462 394 462
use sky130_fd_pr__pfet_01v8_455LYC  sky130_fd_pr__pfet_01v8_455LYC_3
timestamp 1730491634
transform 1 0 -2409 0 1 1123
box -394 -462 394 462
use sky130_fd_pr__pfet_01v8_455LYC  sky130_fd_pr__pfet_01v8_455LYC_4
timestamp 1730491634
transform 1 0 -435 0 1 1123
box -394 -462 394 462
use sky130_fd_pr__pfet_01v8_455LYC  sky130_fd_pr__pfet_01v8_455LYC_5
timestamp 1730491634
transform 1 0 881 0 1 1123
box -394 -462 394 462
<< end >>
