magic
tech sky130A
magscale 1 2
timestamp 1740356695
<< mvpsubdiff >>
rect -161 547 -101 581
rect 4723 547 4783 581
rect -161 521 -127 547
rect -161 -531 -127 -505
rect 4749 521 4783 547
rect 4749 -531 4783 -505
rect -161 -565 -101 -531
rect 4723 -565 4783 -531
<< mvpsubdiffcont >>
rect -101 547 4723 581
rect -161 -505 -127 521
rect 4749 -505 4783 521
rect -101 -565 4723 -531
<< locali >>
rect -506 581 -132 582
rect -506 547 -101 581
rect 4723 547 4783 581
rect -506 521 -127 547
rect -506 -505 -161 521
rect 4749 521 4783 547
rect 470 426 4168 438
rect 470 392 482 426
rect 516 392 566 426
rect 600 392 4034 426
rect 4068 392 4118 426
rect 4152 392 4168 426
rect 470 381 4168 392
rect 470 380 880 381
rect 552 264 880 380
rect 1926 264 2254 381
rect 2384 264 2712 381
rect 3758 380 4168 381
rect 3758 264 4086 380
rect 470 -52 4168 -40
rect 470 -86 482 -52
rect 516 -86 566 -52
rect 600 -86 4034 -52
rect 4068 -86 4118 -52
rect 4152 -86 4168 -52
rect 470 -97 4168 -86
rect 470 -98 880 -97
rect 552 -190 880 -98
rect 1926 -188 2254 -97
rect 2384 -188 2712 -97
rect 3758 -98 4168 -97
rect 3758 -188 4086 -98
rect -506 -531 -127 -505
rect 4749 -531 4783 -505
rect -506 -565 -101 -531
rect 4723 -565 4783 -531
rect -506 -568 -132 -565
<< viali >>
rect 1362 581 1438 582
rect 3200 581 3264 582
rect 4580 581 4628 586
rect -22 547 68 580
rect 1362 547 1438 581
rect 3200 547 3264 581
rect 4580 547 4628 581
rect -22 546 68 547
rect 1362 546 1438 547
rect 3200 546 3264 547
rect 4580 546 4628 547
rect 482 392 516 426
rect 566 392 600 426
rect 4034 392 4068 426
rect 4118 392 4152 426
rect 482 -86 516 -52
rect 566 -86 600 -52
rect 4034 -86 4068 -52
rect 4118 -86 4152 -52
<< metal1 >>
rect -34 580 90 596
rect -34 546 -22 580
rect 68 546 90 580
rect -34 534 90 546
rect 12 304 46 534
rect 470 438 504 640
rect 1350 582 1450 594
rect 1350 546 1362 582
rect 1438 546 1450 582
rect 3188 582 3276 594
rect 3188 546 3200 582
rect 3264 546 3276 582
rect 1350 534 1450 546
rect 1838 540 2008 546
rect 470 426 616 438
rect 470 392 482 426
rect 516 392 566 426
rect 600 392 616 426
rect 470 380 616 392
rect 12 258 140 304
rect 12 210 46 258
rect 12 -148 46 90
rect 470 -40 504 380
rect 1386 298 1420 534
rect 1838 488 1844 540
rect 1896 538 2008 540
rect 1896 488 1950 538
rect 1838 486 1950 488
rect 2002 486 2008 538
rect 1838 482 2008 486
rect 2628 540 2794 546
rect 2628 486 2634 540
rect 2686 488 2730 540
rect 2782 488 2794 540
rect 3188 534 3276 546
rect 2686 486 2794 488
rect 1302 264 1500 298
rect 470 -52 616 -40
rect 470 -86 482 -52
rect 516 -86 566 -52
rect 600 -86 616 -52
rect 470 -98 616 -86
rect 12 -194 126 -148
rect 12 -256 46 -194
rect 470 -250 504 -98
rect 928 -588 962 202
rect 1386 -148 1420 264
rect 1300 -194 1550 -148
rect 1386 -278 1420 -194
rect 1844 -272 1878 482
rect 2628 480 2794 486
rect 2302 -504 2336 224
rect 2760 -268 2794 480
rect 3218 298 3252 534
rect 4134 438 4168 734
rect 4568 586 4640 598
rect 4568 546 4580 586
rect 4628 546 4640 586
rect 4568 534 4640 546
rect 3988 426 4168 438
rect 3988 392 4034 426
rect 4068 392 4118 426
rect 4152 392 4168 426
rect 3988 384 4168 392
rect 4022 380 4168 384
rect 3144 264 3324 298
rect 3218 184 3252 264
rect 3218 -148 3252 96
rect 3128 -194 3378 -148
rect 3218 -270 3252 -194
rect 3676 -236 3710 218
rect 4134 -40 4168 380
rect 4592 304 4626 534
rect 4506 258 4626 304
rect 4592 178 4626 258
rect 3988 -52 4168 -40
rect 3988 -86 4034 -52
rect 4068 -86 4118 -52
rect 4152 -86 4168 -52
rect 3988 -94 4168 -86
rect 4022 -98 4168 -94
rect 4134 -286 4168 -98
rect 4592 -148 4626 62
rect 4500 -194 4626 -148
rect 4592 -250 4626 -194
rect 3676 -588 3710 -398
rect 922 -594 1096 -588
rect 922 -646 928 -594
rect 980 -646 1038 -594
rect 1090 -646 1096 -594
rect 922 -652 1096 -646
rect 3550 -594 3614 -588
rect 3550 -646 3556 -594
rect 3608 -646 3614 -594
rect 3550 -652 3614 -646
rect 3646 -592 3710 -588
rect 3646 -644 3652 -592
rect 3704 -644 3710 -592
rect 3646 -650 3710 -644
<< via1 >>
rect 1844 488 1896 540
rect 1950 486 2002 538
rect 2634 486 2686 540
rect 2730 488 2782 540
rect 928 -646 980 -594
rect 1038 -646 1090 -594
rect 3556 -646 3608 -594
rect 3652 -644 3704 -592
<< metal2 >>
rect 1838 540 2794 546
rect 1838 488 1844 540
rect 1896 538 2634 540
rect 1896 488 1950 538
rect 1838 486 1950 488
rect 2002 486 2634 538
rect 2686 488 2730 540
rect 2782 488 2794 540
rect 2686 486 2794 488
rect 1838 482 2794 486
rect 922 -592 3710 -588
rect 922 -594 3652 -592
rect 922 -646 928 -594
rect 980 -646 1038 -594
rect 1090 -646 3556 -594
rect 3608 -644 3652 -594
rect 3704 -644 3710 -592
rect 3608 -646 3710 -644
rect 922 -650 3710 -646
rect 922 -652 3708 -650
use sky130_fd_pr__nfet_g5v0d10v5_FJPLQ6  sky130_fd_pr__nfet_g5v0d10v5_FJPLQ6_0
timestamp 1740356695
transform 1 0 2319 0 1 -295
box -2319 -157 2319 157
use sky130_fd_pr__nfet_g5v0d10v5_FJPLQ6  sky130_fd_pr__nfet_g5v0d10v5_FJPLQ6_1
timestamp 1740356695
transform 1 0 2319 0 1 157
box -2319 -157 2319 157
<< labels >>
flabel space 170 78 300 150 0 FreeSans 1600 0 0 0 D
flabel space 644 96 774 168 0 FreeSans 800 0 0 0 M10
flabel space 1104 88 1234 160 0 FreeSans 800 0 0 0 D
flabel space 1576 96 1706 168 0 FreeSans 800 0 0 0 D
flabel space 2042 114 2172 186 0 FreeSans 800 0 0 0 M9
flabel space 2476 102 2606 174 0 FreeSans 800 0 0 0 M9
flabel space 2960 96 3090 168 0 FreeSans 800 0 0 0 D
flabel space 3412 92 3542 164 0 FreeSans 800 0 0 0 D
flabel space 3862 106 3992 178 0 FreeSans 800 0 0 0 M10
flabel space 4322 92 4452 164 0 FreeSans 800 0 0 0 D
flabel locali -474 -144 -316 188 0 FreeSans 1600 0 0 0 VSS
port 2 nsew
flabel metal2 2002 482 2634 546 0 FreeSans 1600 0 0 0 IA
port 4 nsew
flabel metal1 470 426 504 640 0 FreeSans 1600 0 0 0 IB
port 5 nsew
flabel metal1 2302 -504 2336 -418 0 FreeSans 1600 0 0 0 IC
port 7 nsew
flabel metal2 1090 -652 3556 -588 0 FreeSans 1600 0 0 0 ID
port 9 nsew
<< end >>
