** sch_path: /foss/designs/OSAD/Learning/Current_mirrors/Design_nmos_current_mirror_ihp_3_3V/simulations/current_mirror_tb_.sch
**.subckt current_mirror_tb_
V1 VDD GND 3.3
V2 VSS GND 0
I0 VDD net2 5u
Vmeas Vout net1 0
.save i(vmeas)
V3 Vout GND 1.65
x1 VSS net2 net1 nmos_current_mirror
**** begin user architecture code

.lib cornerMOShv.lib mos_tt



.param temp=27
.param mm_ok=1
.param mc_ok=1
.control



save all
op
dc V3 0 3.3 0.001
plot i(Vmeas)
wrdata current_mirror.csv i(Vmeas)
.endc


* NGSPICE file created from TOP.ext - technology: ihp-sg13g2

.subckt nmos_current_mirror VSS Iref Iout
X0 VSS Iref Iout VSUB sg13_hv_nmos ad=0.34p pd=2.68u as=0.34p ps=2.68u w=1u l=2.2u
X1 Iout Iref VSS VSUB sg13_hv_nmos ad=0.47302p pd=5.005u as=40.72922p ps=0.14101m w=1u l=2.2u
X2 VSS Iref Iref VSUB sg13_hv_nmos ad=0 pd=0 as=12.88392p ps=59.825u w=1u l=2.2u
X3 Iref VSS VSS VSUB sg13_hv_nmos ad=0 pd=0 as=0 ps=0 w=1u l=2.2u
X4 VSS Iref Iref VSUB sg13_hv_nmos ad=0 pd=0 as=0 ps=0 w=1u l=2.2u
X5 Iref VSS VSS VSUB sg13_hv_nmos ad=0 pd=0 as=0 ps=0 w=1u l=2.2u
X6 VSS Iref Iout VSUB sg13_hv_nmos ad=0 pd=0 as=0 ps=0 w=1u l=2.2u
X7 Iout Iref VSS VSUB sg13_hv_nmos ad=0 pd=0 as=0 ps=0 w=1u l=2.2u
X8 Iref VSS VSS VSUB sg13_hv_nmos ad=0 pd=0 as=0 ps=0 w=1u l=2.2u
X9 VSS Iref Iref VSUB sg13_hv_nmos ad=0 pd=0 as=0 ps=0 w=1u l=2.2u
X10 VSS Iref Iref VSUB sg13_hv_nmos ad=0 pd=0 as=0 ps=0 w=1u l=2.2u
X11 Iref VSS VSS VSUB sg13_hv_nmos ad=0 pd=0 as=0 ps=0 w=1u l=2.2u
C0 VSS Iref 3.04697f
C1 Iref VSUB 5.47165f
C2 VSS VSUB 6.12918f
.ends




**** end user architecture code
**.ends
.GLOBAL GND
.end
