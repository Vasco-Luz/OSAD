** sch_path: /foss/designs/OSAD/Learning/single_ended_amplifiers/Design_and_Analysis_of_Two-Stage_CMOS_Operational_Amplifier_for_Fluorescence_Signal_Processing_sky130_5V/amplifier_design/OTA_AC_TB.sch
**.subckt OTA_AC_TB
V1 VDD GND VDD
V2 VSS GND VSS
Vmeas VDD net2 0
.save i(vmeas)
x5 net2 VSS Va net3 VOUT UUT_VA_sky
C5 VOUT VSS 3p m=1
V16 net1 GND VCM
V17 net3 net1 ac 0.5
V18 net4 VSS ac -0.5
E1 Va net4 net5 VSS 1
R1 VOUT net5 1k ac=1000000000000G m=1
C6 net5 VSS 3p m=1
x6 VDD VSS net8 net7 VOUT_cm UUT_VA_sky
C7 VOUT_cm VSS 3p m=1
V19 net7 net6 VCM
V20 net6 GND ac 1
E2 net8 net6 net9 VSS 1
R2 VOUT_cm net9 1k ac=1000000000000G m=1
C8 net9 VSS 3p m=1
x7 VDD net13 net11 net10 VOUT_a- UUT_VA_sky
C9 VOUT_a- VSS 3p m=1
V21 net10 GND VCM
E3 net11 GND net12 VSS 1
R3 VOUT_a- net12 1k ac=1000000000000G m=1
C10 net12 VSS 3p m=1
V22 net13 VSS ac 1
x8 net14 VSS net16 net15 VOUT_a+ UUT_VA_sky
C11 VOUT_a+ VSS 3p m=1
V23 net15 GND VCM
E4 net16 GND net17 VSS 1
R4 VOUT_a+ net17 1k ac=1000000000000G m=1
C12 net17 VSS 3p m=1
V24 net14 VDD ac 1
x1 VDD VSS net19 VIN+ VOUT_noise UUT_VA_sky
V3 net18 GND VCM
V4 VIN+ net18 ac 0.5
V5 net19 net18 V_OFF
C1 VOUT_noise VSS 3p m=1
**** begin user architecture code
.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice fs

.Temp 27
.param VDD = 5
.param VSS = 0
.param CL = 3p
.param V_OFF = -458.79u
.param VCM=0.9


.control

	save all
	ac dec 100 1 10G
	plot db(v(VOUT)) (180+(180*ph(v(VOUT))/pi))
	plot (db(v(VOUT)) - db(v(VOUT_CM)))
	plot (db(v(VOUT)) - db(v(VOUT_A-)))
	plot (db(v(VOUT))- db(v(VOUT_A+)))
	wrdata VIN_sweep_AC.csv db(v(VOUT)) phase(v(VOUT)) db(v(VOUT_CM)) db(v(VOUT_A-)) db(v(VOUT_A+))

	noise v(VOUT_noise,VSS) V4 dec 10 1 40000k
	print inoise_total
	print onoise_total
	setplot noise1

	plot onoise_spectrum
	plot inoise_spectrum
	op
	print (2.5-V(VOUT))
	print v(VOUT_noise)

.endc




**** end user architecture code
**.ends

* expanding   symbol:  Sky130A/UUT_sky/UUT_VA_sky.sym # of pins=5
** sym_path: /foss/designs/OSAD/LIB/Sky130A/UUT_sky/UUT_VA_sky.sym
** sch_path: /foss/designs/OSAD/LIB/Sky130A/UUT_sky/UUT_VA_sky.sch
.subckt UUT_VA_sky VDD VSS VIN- VIN+ VOUT
*.iopin VDD
*.iopin VSS
*.iopin VIN-
*.iopin VIN+
*.iopin VOUT
x1 VDD VSS VIN+ VIN- VOUT VA001_sky130_1_8V
.ends


* expanding   symbol:  Sky130A/single ended amplifiers/VA001_sky130_1_8V.sym # of pins=5
** sym_path: /foss/designs/OSAD/LIB/Sky130A/single ended amplifiers/VA001_sky130_1_8V.sym
** sch_path: /foss/designs/OSAD/LIB/Sky130A/single ended amplifiers/VA001_sky130_1_8V.sch
.subckt VA001_sky130_1_8V VDD VSS Vin+ Vin- VOUT
*.iopin VDD
*.iopin VSS
*.iopin Vin+
*.iopin Vin-
*.iopin VOUT
XR6 VSS net3 VSS sky130_fd_pr__res_high_po_0p35 L=16 mult=1 m=1
XM1 net1 net2 net3 VSS sky130_fd_pr__nfet_01v8 L=4 W='1 * 8 ' nf=8 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=2
+ m=2
XM2 net2 net2 VSS VSS sky130_fd_pr__nfet_01v8 L=4 W='1 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=2
+ m=2
XM5 VB1 VB1 VDD VDD sky130_fd_pr__pfet_01v8 L=2 W='1 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=2
+ m=2
XM6 VB2 VB1 VDD VDD sky130_fd_pr__pfet_01v8 L=2 W='1 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=2
+ m=2
XM7 net4 VB1 VDD VDD sky130_fd_pr__pfet_01v8 L=2 W='1 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=8
+ m=8
XM10 net5 net5 VSS VSS sky130_fd_pr__nfet_01v8 L=2 W='2.3 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=2
+ m=2
XM11 net6 net5 VSS VSS sky130_fd_pr__nfet_01v8 L=2 W='2.3 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=2
+ m=2
XM12 VOUT VB1 VDD VDD sky130_fd_pr__pfet_01v8 L=2 W='1 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=16
+ m=16
XM14 net7 VB2 net6 VSS sky130_fd_pr__nfet_01v8 L=1.9 W='2 * 1 ' nf=1 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=2
+ m=2
XC1 VOUT net7 sky130_fd_pr__cap_mim_m3_1 W=7.6 L=7.6 MF=4 m=4
XM8 net5 Vin- net4 net4 sky130_fd_pr__pfet_01v8_lvt L=0.8 W='2 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=4
+ m=4
XM9 net6 Vin+ net4 net4 sky130_fd_pr__pfet_01v8_lvt L=0.8 W='2 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=4
+ m=4
XM33 VOUT net6 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.5 W='1.5 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=2
+ m=2
XM3 VB2 VB2 net2 VSS sky130_fd_pr__nfet_01v8_lvt L=2 W='1 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=2
+ m=2
XM4 VB1 VB2 net1 VSS sky130_fd_pr__nfet_01v8_lvt L=2 W='1 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=2
+ m=2
.ends

.GLOBAL GND
.end
