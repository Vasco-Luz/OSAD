magic
tech sky130A
magscale 1 2
timestamp 1738953643
<< nwell >>
rect -394 -214 394 248
<< pmos >>
rect -300 -114 300 186
<< pdiff >>
rect -358 174 -300 186
rect -358 -102 -346 174
rect -312 -102 -300 174
rect -358 -114 -300 -102
rect 300 174 358 186
rect 300 -102 312 174
rect 346 -102 358 174
rect 300 -114 358 -102
<< pdiffc >>
rect -346 -102 -312 174
rect 312 -102 346 174
<< poly >>
rect -300 186 300 212
rect -300 -161 300 -114
rect -300 -178 -227 -161
rect -243 -195 -227 -178
rect 227 -178 300 -161
rect 227 -195 243 -178
rect -243 -211 243 -195
<< polycont >>
rect -227 -195 227 -161
<< locali >>
rect -346 174 -312 190
rect -346 -118 -312 -102
rect 312 174 346 190
rect 312 -118 346 -102
rect -243 -195 -227 -161
rect 227 -195 243 -161
<< viali >>
rect -346 -102 -312 174
rect 312 -102 346 174
rect -227 -195 227 -161
<< metal1 >>
rect -352 174 -306 516
rect -352 -102 -346 174
rect -312 -102 -306 174
rect -352 -114 -306 -102
rect 306 174 352 330
rect 306 -102 312 174
rect 346 -102 352 174
rect 306 -114 352 -102
rect -346 -132 -312 -114
rect -239 -161 239 -155
rect -239 -195 -227 -161
rect 227 -195 239 -161
rect -239 -201 239 -195
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.5 l 3 m 1 nf 1 diffcov 100 polycov 80 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 80 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
