** sch_path:
*+ /home/vasco/Desktop/sky130A/amplifiers/single_stage_amps/basic_stages/cs_resistor_stage/full_script/cs_resistor_stage_test.sch
**.subckt cs_resistor_stage_test
Vmeas VDD net1 0
.save i(vmeas)
V1 VDD GND 5
.save i(v1)
V2 VIN GND 1.265
.save i(v2)
V3 VINT GND ac 1.0 sin (0 100u 100k)
.save i(v3)
R2 VOUT GND 10G m=1
C1 VINT net2 1 m=1
R3 VIN net2 10M m=1
R5 VOUTT GND 10G m=1
XM1 VOUT VIN GND GND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=60 nf=10 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
C2 net3 VOUTT 100u m=1
XR6 VOUT net1 VDD sky130_fd_pr__res_high_po_0p35 L=1*8 mult=2 m=2
x1 VDD GND net2 net3 cs_resistor_stage
**** begin user architecture code

**************************************************************
**************************************************************
**************************************************************
**************************************************************
**************************************************************
*LIBs*********************************************************
**************************************************************
**************************************************************
**************************************************************
**************************************************************
**************************************************************
*.lib /home/vasco/Desktop/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
* chose the corners in the corner file
* tt_mm for mismatch
* ss ff sf fs standart corners
* ll hh lh hl capacitor and resistors corners
* mc for total process variation including corners
**************************************************************
**************************************************************
**************************************************************
**************************************************************
**************************************************************
*Corners/montecarlo options***********************************
**************************************************************
**************************************************************
**************************************************************
**************************************************************
**************************************************************
.TEMP 27
**************************************************************
**************************************************************
**************************************************************
**************************************************************
*SIMULATION and Plots*****************************************
**************************************************************
**************************************************************
**************************************************************
**************************************************************
.control
save all
dc V2 0 3.3 0.01
*dc simulation
plot v(VOUT) v(VIN) deriv(v(VOUT))
*ploting VIN VOUT and the voltage gain
plot i(Vmeas)
*ploting the current for curiosity
tran 0.1ns 20u
*transient simulation
plot (v(VINT)) (v(VOUTT))
*simple plot to exemplify the gain
fft v(VOUTT) v(VINT)
*fast fourier transfor
plot mag(v(VOUTT)) mag(v(VINT))
* analyse the frequency spectrum of the transient waves, to detect distortion
ac dec 20 1 50G
*simple ac simulation
plot v(VOUTT) v(VOUTT)
*gain in function of the input frequency
.endc


.param mc_mm_switch=0
.param mc_pr_switch=0
.include /home/vasco/Desktop/pdk/sky130A/libs.tech/ngspice/corners/tt.spice
.include /home/vasco/Desktop/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/vasco/Desktop/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/vasco/Desktop/pdk/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends

* expanding   symbol:
*+  /home/vasco/Desktop/sky130A/amplifiers/single_stage_amps/basic_stages/cs_resistor_stage/cs_resistor_stage.sym # of pins=4
** sym_path:
*+ /home/vasco/Desktop/sky130A/amplifiers/single_stage_amps/basic_stages/cs_resistor_stage/cs_resistor_stage.sym
** sch_path:
*+ /home/vasco/Desktop/sky130A/amplifiers/single_stage_amps/basic_stages/cs_resistor_stage/cs_resistor_stage.sch
.subckt cs_resistor_stage VDD VSS VIN VOUT
*.iopin VDD
*.iopin VSS
*.iopin VIN
*.iopin VOUT
XM1 VOUT VIN VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=60 nf=10 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XR6 VOUT VDD VDD sky130_fd_pr__res_high_po_0p35 L=1*8 mult=2 m=2
.ends

.GLOBAL GND
.end
