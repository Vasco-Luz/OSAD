magic
tech sky130A
magscale 1 2
timestamp 1730506627
<< locali >>
rect 10 2554 4410 2560
rect 10 2520 20 2554
rect 4398 2520 4410 2554
rect 10 2510 4410 2520
rect 250 1412 304 2510
rect 250 1328 762 1412
rect 250 350 304 1328
rect 248 250 304 350
rect 1566 304 1620 2510
rect 2882 326 2936 2510
rect 4194 1414 4248 2510
rect 3744 1326 4248 1414
rect 4194 250 4248 1326
rect 248 166 760 250
rect 3746 160 4248 250
<< viali >>
rect 20 2520 4398 2554
<< metal1 >>
rect -16 2554 4420 2570
rect -16 2520 20 2554
rect 4398 2520 4420 2554
rect -16 2500 4420 2520
rect 910 1480 958 2312
rect 911 1284 957 1480
rect 894 1230 904 1284
rect 964 1230 974 1284
rect 911 132 957 1230
rect 888 80 898 132
rect 970 80 980 132
rect 911 -99 957 80
rect 2226 -36 2274 2310
rect 3542 1284 3590 2310
rect 3526 1228 3536 1284
rect 3594 1228 3604 1284
rect 3542 132 3590 1228
rect 3518 78 3528 132
rect 3604 78 3614 132
rect 3542 -48 3590 78
<< via1 >>
rect 904 1230 964 1284
rect 898 80 970 132
rect 3536 1228 3594 1284
rect 3528 78 3604 132
<< metal2 >>
rect 904 1284 964 1294
rect 1132 1270 1192 1372
rect 1790 1270 1850 1374
rect 2658 1270 2718 1374
rect 3316 1270 3376 1370
rect 3536 1284 3594 1294
rect 964 1240 3536 1270
rect 904 1220 964 1230
rect 3536 1218 3594 1228
rect 898 132 970 142
rect 1132 120 1192 220
rect 1790 120 1850 222
rect 2658 120 2718 214
rect 3316 120 3376 220
rect 3528 132 3604 142
rect 970 88 3528 120
rect 898 70 970 80
rect 3528 68 3604 78
use PMOS_cell  PMOS_cell_0 ~/Desktop/OSAD/my_ip/Layouts/VA001_PMOS_1.8_sky130
timestamp 1730503605
transform 1 0 211 0 1 157
box -227 -161 4223 2431
<< labels >>
flabel space 466 1788 752 2110 0 FreeSans 800 0 0 0 Dummy
flabel space 494 716 780 1038 0 FreeSans 800 0 0 0 Dummy
flabel space 3746 592 4032 914 0 FreeSans 800 0 0 0 Dummy
flabel space 3722 1730 4008 2052 0 FreeSans 800 0 0 0 Dummy
flabel space 1146 1782 1400 2160 0 FreeSans 800 0 0 0 M1
flabel space 1106 620 1360 998 0 FreeSans 800 0 0 0 M1
flabel space 3046 592 3300 970 0 FreeSans 800 0 0 0 M1
flabel space 3684 1018 3938 1396 0 FreeSans 800 0 0 0 M1
flabel space 1814 648 2044 922 0 FreeSans 800 0 0 0 M2
flabel space 2464 604 2694 878 0 FreeSans 800 0 0 0 M2
flabel space 2442 1772 2672 2046 0 FreeSans 800 0 0 0 M2
flabel space 1848 1758 2078 2032 0 FreeSans 800 0 0 0 M2
<< end >>
