* NGSPICE file created from Nmos_lower_current_mirror.ext - technology: sky130A

.subckt Nmos_lower_current_mirror VSS IC ID IE 
X0 IC VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3.2
X1 ID VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.16003 pd=10.325 as=2.32002 ps=20.645 w=1 l=3.2
X2 IC VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=2.90002 pd=25.805 as=0 ps=0 w=1 l=3.2
X3 ID VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=3.2
X4 ID VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=3.2
X5 VSS ID ID VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3.2
X6 IC VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=3.2
X7 VSS ID ID VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=3.2
X8 ID VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=3.2
X9 IC VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=3.2
X10 IE ID IC VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=3.2
X11 IC ID IE VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=3.2
X12 VSS ID ID VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=3.2
X13 VSS ID ID VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=3.2
X14 IE ID IC VSS sky130_fd_pr__nfet_g5v0d10v5 ad=2.32 pd=20.64 as=0 ps=0 w=1 l=3.2
X15 IC ID IE VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=3.2
X16 IE ID IC VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=3.2
X17 IC ID IE VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=3.2
X18 IE ID IC VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=3.2
X19 IC ID IE VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=3.2
X20 IE ID IC VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=3.2
X21 IC ID IE VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=3.2
X22 IE ID IC VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=3.2
X23 IC ID IE VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=3.2
X24 IE ID IC VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=3.2
X25 IC ID IE VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=3.2
X26 IE ID IC VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=3.2
X27 IC ID IE VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=3.2
C0 IE IC 3.21167f
C1 ID IC 2.55348f
C2 VSS ID 6.7579f
C3 IE 0 2.10306f
C4 ID 0 21.8586f
C5 VSS 0 2.30348f
C6 IC 0 2.30032f
.ends
