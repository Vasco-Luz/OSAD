** sch_path: /foss/pdks/ihp-sg13g2/libs.tech/xschem/sg13g2_tests/mc_mim_cap_ac.sch
**.subckt mc_mim_cap_ac
V1 in GND dc 0 ac 1
R2 out GND 100k m=1
XC1 out in cap_cmim w=7.0e-6 l=7.0e-6 m=1
**** begin user architecture code


.param mc_ok = 1
.control
let mc_runs = 1000
let run = 0
shell rm mc_cmim.csv
***************** LOOP *********************
dowhile run < mc_runs
reset
set run=$&run
save all
ac dec 1000 1e6 100e9
let mag=abs(out)
meas ac freq_at when mag = 0.707
let C = 1/(2*PI*freq_at*1e+5)
print C >> mc_cmim.csv
let run=run+1
end
***************** LOOP *********************
.endc



.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerCAP.lib cap_wcs_stat

**** end user architecture code
**.ends
.GLOBAL GND
.end
