* NGSPICE file created from pmos_current_mirror.ext - technology: sky130A

.subckt pmos_current_mirror VDD IB IA
X0 IA IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=3
X1 IA IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=14.3 as=1.74 ps=14.3 w=1.5 l=3
X2 IA IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1.5 l=3
X3 IA IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1.5 l=3
X4 VDD IA IB VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.218 ps=1.79 w=1.5 l=3
X5 IB IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.218 pd=1.79 as=0.435 ps=3.58 w=1.5 l=3
X6 VDD IA IB VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.87 ps=7.16 w=1.5 l=3
X7 IB IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1.5 l=3
C0 VDD IA 6.5f
C1 VDD VSUBS 14.6f
C2 IA VSUBS 3.95f
.ends
