** sch_path: /foss/designs/OSAD/Learning/single_ended_amplifiers/A_High_Precision_Micropower_Operational_Amplifier_IHP130_3_3/current_reference/testbench.sch
**.subckt testbench
VDD VDD GND 5
VSS VSS GND 0
XR2 net1 Va rppd w=0.5e-6 l=5e-6 m=1 b=0
XQ1 net1 Va VSS VSS npn13G2v Nx=1
Vmeas net4 net5 0
.save i(vmeas)
XM1 net2 net2 VDD VDD sg13_hv_pmos w=1.0u l=4u ng=1 m=2
XM2 Va Va net2 net2 sg13_hv_pmos w=1.0u l=4u ng=1 m=2
XQ2 net4 net3 VDD pnpMPA a=2e-12 p=6e-06 m=1
XQ3 net5 net1 VSS VSS npn13G2v Nx=2
XQ4 VSS net4 net3 pnpMPA a=2e-12 p=6e-06 m=1
**** begin user architecture code

.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerHBT.lib hbt_typ


.lib cornerMOShv.lib mos_tt


.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerRES.lib res_typ_stat



.param temp=27
.param mm_ok=1
.param mc_ok=1
.control
save all
dc temp -40 125 1
plot i(Vmeas)
plot v(Va)
dc VDD 3 6 0.01
plot i(Vmeas)
plot v(Va)
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
