magic
tech sky130A
magscale 1 2
timestamp 1740408217
<< error_p >>
rect -574 -198 -544 130
rect -508 -132 -478 64
rect 478 -132 508 64
rect -508 -136 508 -132
rect 544 -198 574 130
rect -574 -202 574 -198
<< nwell >>
rect -544 -198 544 164
<< mvpmos >>
rect -450 -136 450 64
<< mvpdiff >>
rect -508 52 -450 64
rect -508 -124 -496 52
rect -462 -124 -450 52
rect -508 -136 -450 -124
rect 450 52 508 64
rect 450 -124 462 52
rect 496 -124 508 52
rect 450 -136 508 -124
<< mvpdiffc >>
rect -496 -124 -462 52
rect 462 -124 496 52
<< poly >>
rect -363 145 363 161
rect -363 128 -347 145
rect -450 111 -347 128
rect 347 128 363 145
rect 347 111 450 128
rect -450 64 450 111
rect -450 -162 450 -136
<< polycont >>
rect -347 111 347 145
<< locali >>
rect -363 111 -347 145
rect 347 111 363 145
rect -496 52 -462 68
rect -496 -140 -462 -124
rect 462 52 496 68
rect 462 -140 496 -124
<< viali >>
rect -347 111 347 145
rect -496 -124 -462 52
rect 462 -124 496 52
<< metal1 >>
rect -359 145 359 151
rect -359 111 -347 145
rect 347 111 359 145
rect -359 105 359 111
rect -502 52 -456 64
rect -502 -124 -496 52
rect -462 -124 -456 52
rect -502 -136 -456 -124
rect 456 52 502 64
rect 456 -124 462 52
rect 496 -124 502 52
rect 456 -136 502 -124
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1 l 4.5 m 1 nf 1 diffcov 100 polycov 80 guard 0 glc 0 grc 0 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 80 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
