magic
tech sky130A
magscale 1 2
timestamp 1693785227
<< locali >>
rect -312 3674 -260 3834
rect 1182 3680 1234 3840
<< viali >>
rect 3150 6470 3190 6550
rect 3100 1504 3140 1584
<< metal1 >>
rect 3120 6550 3220 6622
rect 3120 6470 3150 6550
rect 3190 6470 3220 6550
rect 3120 6392 3220 6470
rect 2980 6344 3362 6392
rect 2980 5388 3362 5440
rect 3120 5356 3220 5388
rect 3120 5304 3134 5356
rect 3208 5304 3220 5356
rect 3120 5294 3220 5304
rect -643 3922 -92 3980
rect -314 3288 -258 3812
rect -150 3764 -92 3922
rect 1016 3890 2492 3942
rect 20 3812 236 3814
rect 352 3812 568 3814
rect 684 3812 904 3814
rect -148 3288 -92 3764
rect 18 3772 240 3812
rect 18 3288 74 3772
rect 184 3288 240 3772
rect 350 3772 572 3812
rect 350 3288 406 3772
rect 516 3288 572 3772
rect 682 3772 904 3812
rect 682 3302 740 3772
rect 682 3288 738 3302
rect 848 3290 904 3772
rect 1016 3290 1068 3890
rect 3076 3864 3248 3870
rect 3076 3800 3082 3864
rect 3242 3800 3248 3864
rect 3076 3794 3248 3800
rect -146 2610 -90 3092
rect 18 2610 74 3092
rect -146 2568 74 2610
rect 186 2610 242 3092
rect 348 2610 404 3092
rect 186 2568 404 2610
rect 516 2610 572 3092
rect 684 2610 740 3092
rect 516 2568 740 2610
rect 848 2610 904 3090
rect 1014 2610 1070 3092
rect 848 2566 1070 2610
rect 3070 1584 3180 1590
rect 3070 1512 3100 1584
rect 3140 1512 3180 1584
rect 3070 1460 3090 1512
rect 3160 1460 3180 1512
rect 3070 1450 3180 1460
rect 2934 1394 3318 1450
rect 2934 438 3318 498
rect 3080 140 3162 438
<< via1 >>
rect 3134 5304 3208 5356
rect 3082 3800 3242 3864
rect 3132 3356 3196 3470
rect 3090 1504 3100 1512
rect 3100 1504 3140 1512
rect 3140 1504 3160 1512
rect 3090 1460 3160 1504
<< metal2 >>
rect 3128 5356 3214 5362
rect 3128 5304 3134 5356
rect 3208 5304 3214 5356
rect 3128 3870 3214 5304
rect 3076 3864 3248 3870
rect 3076 3800 3082 3864
rect 3242 3800 3248 3864
rect 3076 3794 3248 3800
rect 3084 3470 3202 3476
rect 3084 3356 3132 3470
rect 3196 3356 3202 3470
rect 3084 3330 3202 3356
rect 3084 1512 3166 3330
rect 3084 1460 3090 1512
rect 3160 1460 3166 1512
rect 3084 1454 3166 1460
use sky130_fd_pr__res_high_po_0p35_G4FHUE  sky130_fd_pr__res_high_po_0p35_G4FHUE_0
timestamp 1693784648
transform 1 0 3126 0 1 957
box -428 -657 428 657
use sky130_fd_pr__res_high_po_0p35_G4FHUE  sky130_fd_pr__res_high_po_0p35_G4FHUE_1
timestamp 1693784648
transform 1 0 3170 0 1 5903
box -428 -657 428 657
use sky130_fd_pr__res_high_po_0p35_XKGYDU  sky130_fd_pr__res_high_po_0p35_XKGYDU_0
timestamp 1693784648
transform -1 0 461 0 -1 3185
box -1009 -707 1009 707
use sky130_fd_pr__rf_npn_05v5_W1p00L2p00  sky130_fd_pr__rf_npn_05v5_W1p00L2p00_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1692646696
transform 1 0 2304 0 1 2468
box 0 0 1724 1924
<< labels >>
flabel metal1 -643 3922 -92 3980 0 FreeSans 1600 0 0 0 VDD
port 1 nsew
flabel metal1 3080 140 3162 498 0 FreeSans 1600 0 0 0 VSS
port 3 nsew
flabel metal1 3120 6550 3220 6622 0 FreeSans 1600 0 0 0 VIN
port 5 nsew
flabel metal2 3128 3864 3214 5304 0 FreeSans 1600 0 0 0 VOUT
port 7 nsew
<< end >>
