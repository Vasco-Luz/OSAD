* NGSPICE file created from cs_current_pmos_stage_post.ext - technology: sky130A

.subckt cs_current_pmos_stage_post VDD VSS VIN VOUT VB
X0 VOUT VB VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.8
X1 VDD VB VOUT VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.8
X2 VOUT VB VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.8
X3 VDD VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.8
X4 VDD VB VOUT VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.8
X5 VOUT VB VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.8
X6 VDD VB VOUT VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.8
X7 VOUT VB VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.8
X8 VDD VB VOUT VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.8
X9 VOUT VB VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.8
X10 VDD VB VOUT VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.8
X11 VDD VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.8
X12 VSS VSS VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=2.32 pd=16.6 as=1.16 ps=8.29 w=8 l=0.8
X13 VSS VIN VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.8
X14 VOUT VIN VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.8
X15 VSS VIN VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.8
X16 VOUT VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=2.32 ps=16.6 w=8 l=0.8
X17 VOUT VIN VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.8
X18 VSS VIN VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.8
X19 VOUT VIN VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.8
X20 VOUT VIN VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.8
X21 VSS VIN VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.8
X22 VSS VIN VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.8
X23 VOUT VIN VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.8
C0 VOUT VIN 2.97f
C1 VOUT VSS 6.95f
C2 VSS VIN 2.08f
C3 VDD VB 4.45f
C4 VOUT VDD 3.31f
C5 VSS 0 3.49f
C6 VIN 0 3.13f
C7 VOUT 0 2.07f
C8 VDD 0 14.6f
.ends
