magic
tech sky130A
magscale 1 2
timestamp 1740347700
<< error_p >>
rect -1091 -198 -1061 130
rect -1025 -132 -995 64
rect 995 -132 1025 64
rect -1025 -136 1025 -132
rect 1061 -198 1091 130
rect -1091 -202 1091 -198
<< nwell >>
rect -1061 -198 1061 164
<< mvpmos >>
rect -967 -136 -527 64
rect -469 -136 -29 64
rect 29 -136 469 64
rect 527 -136 967 64
<< mvpdiff >>
rect -1025 52 -967 64
rect -1025 -124 -1013 52
rect -979 -124 -967 52
rect -1025 -136 -967 -124
rect -527 52 -469 64
rect -527 -124 -515 52
rect -481 -124 -469 52
rect -527 -136 -469 -124
rect -29 52 29 64
rect -29 -124 -17 52
rect 17 -124 29 52
rect -29 -136 29 -124
rect 469 52 527 64
rect 469 -124 481 52
rect 515 -124 527 52
rect 469 -136 527 -124
rect 967 52 1025 64
rect 967 -124 979 52
rect 1013 -124 1025 52
rect 967 -136 1025 -124
<< mvpdiffc >>
rect -1013 -124 -979 52
rect -515 -124 -481 52
rect -17 -124 17 52
rect 481 -124 515 52
rect 979 -124 1013 52
<< poly >>
rect -926 145 -568 161
rect -926 128 -910 145
rect -967 111 -910 128
rect -584 128 -568 145
rect -428 145 -70 161
rect -428 128 -412 145
rect -584 111 -527 128
rect -967 64 -527 111
rect -469 111 -412 128
rect -86 128 -70 145
rect 70 145 428 161
rect 70 128 86 145
rect -86 111 -29 128
rect -469 64 -29 111
rect 29 111 86 128
rect 412 128 428 145
rect 568 145 926 161
rect 568 128 584 145
rect 412 111 469 128
rect 29 64 469 111
rect 527 111 584 128
rect 910 128 926 145
rect 910 111 967 128
rect 527 64 967 111
rect -967 -162 -527 -136
rect -469 -162 -29 -136
rect 29 -162 469 -136
rect 527 -162 967 -136
<< polycont >>
rect -910 111 -584 145
rect -412 111 -86 145
rect 86 111 412 145
rect 584 111 910 145
<< locali >>
rect -926 111 -910 145
rect -584 111 -568 145
rect -428 111 -412 145
rect -86 111 -70 145
rect 70 111 86 145
rect 412 111 428 145
rect 568 111 584 145
rect 910 111 926 145
rect -1013 52 -979 68
rect -1013 -140 -979 -124
rect -515 52 -481 68
rect -515 -140 -481 -124
rect -17 52 17 68
rect -17 -140 17 -124
rect 481 52 515 68
rect 481 -140 515 -124
rect 979 52 1013 68
rect 979 -140 1013 -124
<< viali >>
rect -910 111 -584 145
rect -412 111 -86 145
rect 86 111 412 145
rect 584 111 910 145
rect -1013 -124 -979 52
rect -515 -124 -481 52
rect -17 -124 17 52
rect 481 -124 515 52
rect 979 -124 1013 52
<< metal1 >>
rect -922 145 -572 151
rect -922 111 -910 145
rect -584 111 -572 145
rect -922 105 -572 111
rect -424 145 -74 151
rect -424 111 -412 145
rect -86 111 -74 145
rect -424 105 -74 111
rect 74 145 424 151
rect 74 111 86 145
rect 412 111 424 145
rect 74 105 424 111
rect 572 145 922 151
rect 572 111 584 145
rect 910 111 922 145
rect 572 105 922 111
rect -1019 52 -973 64
rect -1019 -124 -1013 52
rect -979 -124 -973 52
rect -1019 -136 -973 -124
rect -521 52 -475 64
rect -521 -124 -515 52
rect -481 -124 -475 52
rect -521 -136 -475 -124
rect -23 52 23 64
rect -23 -124 -17 52
rect 17 -124 23 52
rect -23 -136 23 -124
rect 475 52 521 64
rect 475 -124 481 52
rect 515 -124 521 52
rect 475 -136 521 -124
rect 973 52 1019 64
rect 973 -124 979 52
rect 1013 -124 1019 52
rect 973 -136 1019 -124
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1 l 2.2 m 1 nf 4 diffcov 100 polycov 80 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 80 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
