* NGSPICE file created from VA001_sky130_5V.ext - technology: sky130A

.subckt VA001_sky130_5V VDD VSS Vin+ Vin- VOUT
X0 bias_res_0/li_3975_7364# Lower_Nmos_0/IC VSS sky130_fd_pr__res_xhigh_po_0p69 l=1.62
X1 bias_res_0/li_5098_7502# bias_res_0/li_3975_7364# VSS sky130_fd_pr__res_xhigh_po_0p69 l=1.62
X2 VSS bias_res_0/res_poly$1_2/a_n69_n582# VSS sky130_fd_pr__res_xhigh_po_0p69 l=1.62
X3 VSS bias_res_0/res_poly$1_3/a_n69_n582# VSS sky130_fd_pr__res_xhigh_po_0p69 l=1.62
X4 bias_res_0/li_5098_7502# bias_res_0/li_3975_7618# VSS sky130_fd_pr__res_xhigh_po_0p69 l=1.62
X5 bias_res_0/li_5098_8010# bias_res_0/li_3974_7872# VSS sky130_fd_pr__res_xhigh_po_0p69 l=1.62
X6 bias_res_0/li_5098_8010# bias_res_0/li_3975_8126# VSS sky130_fd_pr__res_xhigh_po_0p69 l=1.62
X7 VSS bias_res_0/li_3975_8380# VSS sky130_fd_pr__res_xhigh_po_0p69 l=1.62
X8 bias_res_0/li_3975_7618# bias_res_0/li_2811_7755# VSS sky130_fd_pr__res_xhigh_po_0p69 l=1.62
X9 bias_res_0/res_poly$1_9/a_n69_146# VSS VSS sky130_fd_pr__res_xhigh_po_0p69 l=1.62
X10 bias_res_0/li_3974_7872# bias_res_0/li_2811_7755# VSS sky130_fd_pr__res_xhigh_po_0p69 l=1.62
X11 bias_res_0/res_poly$1_11/a_n69_146# VSS VSS sky130_fd_pr__res_xhigh_po_0p69 l=1.62
X12 bias_res_0/li_3975_8126# bias_res_0/li_2811_8263# VSS sky130_fd_pr__res_xhigh_po_0p69 l=1.62
X13 bias_res_0/li_3975_8380# bias_res_0/li_2811_8263# VSS sky130_fd_pr__res_xhigh_po_0p69 l=1.62
X14 VOUT VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1 pd=4.5 as=1.2 ps=8.6 w=4 l=1
X15 VSS active_load_0/IA VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1 pd=4.5 as=1 ps=4.5 w=4 l=1
X16 VSS VSS VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.2 pd=8.6 as=1 ps=4.5 w=4 l=1
X17 VOUT active_load_0/IA VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1 pd=4.5 as=1 ps=4.5 w=4 l=1
X18 VOUT VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=8 pd=36 as=20 ps=127.6 w=4 l=1
X19 VSS active_load_0/IA VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4 l=1
X20 VSS VSS VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4 l=1
X21 VOUT active_load_0/IA VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4 l=1
X22 VSS active_load_0/IB active_load_0/IA VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.375 pd=2 as=0.375 ps=2 w=1.5 l=2
X23 active_load_0/IB VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.375 pd=2 as=0.45 ps=3.6 w=1.5 l=2
X24 active_load_0/IA active_load_0/IB VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.375 pd=2 as=0.375 ps=2 w=1.5 l=2
X25 VSS active_load_0/IB active_load_0/IB VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.375 pd=2 as=0.375 ps=2 w=1.5 l=2
X26 VSS VSS active_load_0/IB VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.45 pd=3.6 as=0.375 ps=2 w=1.5 l=2
X27 active_load_0/IB active_load_0/IB VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.375 pd=2 as=0.375 ps=2 w=1.5 l=2
X28 VSS active_load_0/IB active_load_0/IA VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=2.34 ps=14.8 w=1.5 l=2
X29 active_load_0/IB VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=3 pd=16 as=0 ps=0 w=1.5 l=2
X30 active_load_0/IA active_load_0/IB VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1.5 l=2
X31 VSS active_load_0/IB active_load_0/IB VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1.5 l=2
X32 VSS VSS active_load_0/IB VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1.5 l=2
X33 active_load_0/IB active_load_0/IB VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1.5 l=2
X34 active_load_0/IA Vin+ Pmos_current_mirror_0/IC Pmos_current_mirror_0/IC sky130_fd_pr__pfet_g5v0d10v5 ad=1.125 pd=5 as=1.125 ps=5 w=4.5 l=1
X35 active_load_0/IB Vin- Pmos_current_mirror_0/IC Pmos_current_mirror_0/IC sky130_fd_pr__pfet_g5v0d10v5 ad=1.125 pd=5 as=1.125 ps=5 w=4.5 l=1
X36 Pmos_current_mirror_0/IC Pmos_current_mirror_0/IC Pmos_current_mirror_0/IC Pmos_current_mirror_0/IC sky130_fd_pr__pfet_g5v0d10v5 ad=1.125 pd=5 as=1.35 ps=9.6 w=4.5 l=1
X37 Pmos_current_mirror_0/IC Pmos_current_mirror_0/IC Pmos_current_mirror_0/IC Pmos_current_mirror_0/IC sky130_fd_pr__pfet_g5v0d10v5 ad=1.35 pd=9.6 as=1.125 ps=5 w=4.5 l=1
X38 active_load_0/IB Vin- Pmos_current_mirror_0/IC Pmos_current_mirror_0/IC sky130_fd_pr__pfet_g5v0d10v5 ad=1.125 pd=5 as=1.125 ps=5 w=4.5 l=1
X39 active_load_0/IA Vin+ Pmos_current_mirror_0/IC Pmos_current_mirror_0/IC sky130_fd_pr__pfet_g5v0d10v5 ad=1.125 pd=5 as=1.125 ps=5 w=4.5 l=1
X40 Pmos_current_mirror_0/IC Vin+ active_load_0/IA Pmos_current_mirror_0/IC sky130_fd_pr__pfet_g5v0d10v5 ad=1.125 pd=5 as=1.125 ps=5 w=4.5 l=1
X41 Pmos_current_mirror_0/IC Vin+ active_load_0/IA Pmos_current_mirror_0/IC sky130_fd_pr__pfet_g5v0d10v5 ad=1.125 pd=5 as=1.125 ps=5 w=4.5 l=1
X42 Pmos_current_mirror_0/IC Vin- active_load_0/IB Pmos_current_mirror_0/IC sky130_fd_pr__pfet_g5v0d10v5 ad=1.125 pd=5 as=1.125 ps=5 w=4.5 l=1
X43 Pmos_current_mirror_0/IC Vin- active_load_0/IB Pmos_current_mirror_0/IC sky130_fd_pr__pfet_g5v0d10v5 ad=1.125 pd=5 as=1.125 ps=5 w=4.5 l=1
X44 active_load_0/IB Vin- Pmos_current_mirror_0/IC Pmos_current_mirror_0/IC sky130_fd_pr__pfet_g5v0d10v5 ad=9 pd=40 as=31.9 ps=162.39999 w=4.5 l=1
X45 active_load_0/IA Vin+ Pmos_current_mirror_0/IC Pmos_current_mirror_0/IC sky130_fd_pr__pfet_g5v0d10v5 ad=9 pd=40 as=0 ps=0 w=4.5 l=1
X46 Pmos_current_mirror_0/IC Pmos_current_mirror_0/IC Pmos_current_mirror_0/IC Pmos_current_mirror_0/IC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4.5 l=1
X47 Pmos_current_mirror_0/IC Pmos_current_mirror_0/IC Pmos_current_mirror_0/IC Pmos_current_mirror_0/IC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4.5 l=1
X48 active_load_0/IA Vin+ Pmos_current_mirror_0/IC Pmos_current_mirror_0/IC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4.5 l=1
X49 active_load_0/IB Vin- Pmos_current_mirror_0/IC Pmos_current_mirror_0/IC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4.5 l=1
X50 Pmos_current_mirror_0/IC Vin- active_load_0/IB Pmos_current_mirror_0/IC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4.5 l=1
X51 Pmos_current_mirror_0/IC Vin- active_load_0/IB Pmos_current_mirror_0/IC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4.5 l=1
X52 Pmos_current_mirror_0/IC Vin+ active_load_0/IA Pmos_current_mirror_0/IC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4.5 l=1
X53 Pmos_current_mirror_0/IC Vin+ active_load_0/IA Pmos_current_mirror_0/IC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4.5 l=1
X54 VDD Pmos_current_mirror_0/IA Pmos_current_mirror_0/IA VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2.2
X55 VDD Pmos_current_mirror_0/IA VOUT VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2.2
X56 Pmos_current_mirror_0/IA VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.3 ps=2.6 w=1 l=2.2
X57 VOUT Pmos_current_mirror_0/IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2.2
X58 Pmos_current_mirror_0/IC Pmos_current_mirror_0/IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2.2
X59 VDD Pmos_current_mirror_0/IA Pmos_current_mirror_0/IB VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2.2
X60 VDD VDD Pmos_current_mirror_0/IA VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2.2
X61 VDD Pmos_current_mirror_0/IA Pmos_current_mirror_0/IC VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2.2
X62 VDD Pmos_current_mirror_0/IA Pmos_current_mirror_0/IC VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2.2
X63 VOUT Pmos_current_mirror_0/IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2.2
X64 VOUT Pmos_current_mirror_0/IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2.2
X65 VOUT Pmos_current_mirror_0/IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2.2
X66 Pmos_current_mirror_0/IB Pmos_current_mirror_0/IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2.2
X67 Pmos_current_mirror_0/IA Pmos_current_mirror_0/IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2.2
X68 Pmos_current_mirror_0/IC Pmos_current_mirror_0/IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2.2
X69 VDD Pmos_current_mirror_0/IA VOUT VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2.2
X70 VDD Pmos_current_mirror_0/IA VOUT VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2.2
X71 VDD Pmos_current_mirror_0/IA VOUT VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2.2
X72 VDD Pmos_current_mirror_0/IA VOUT VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2.2
X73 VDD Pmos_current_mirror_0/IA VOUT VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2.2
X74 Pmos_current_mirror_0/IC Pmos_current_mirror_0/IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2.2
X75 VDD VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.3 pd=2.6 as=0.25 ps=1.5 w=1 l=2.2
X76 Pmos_current_mirror_0/IC Pmos_current_mirror_0/IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2.2
X77 VOUT Pmos_current_mirror_0/IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2.2
X78 VOUT Pmos_current_mirror_0/IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2.2
X79 VOUT Pmos_current_mirror_0/IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2.2
X80 VOUT Pmos_current_mirror_0/IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2.2
X81 VDD Pmos_current_mirror_0/IA VOUT VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2.2
X82 VDD Pmos_current_mirror_0/IA VOUT VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2.2
X83 VDD Pmos_current_mirror_0/IA Pmos_current_mirror_0/IC VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2.2
X84 VDD Pmos_current_mirror_0/IA Pmos_current_mirror_0/IC VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2.2
X85 VDD Pmos_current_mirror_0/IA Pmos_current_mirror_0/IA VDD sky130_fd_pr__pfet_g5v0d10v5 ad=16.2 pd=100.4 as=2 ps=12 w=1 l=2.2
X86 VDD Pmos_current_mirror_0/IA VOUT VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=8 ps=48 w=1 l=2.2
X87 Pmos_current_mirror_0/IA VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=2.2
X88 VOUT Pmos_current_mirror_0/IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=2.2
X89 Pmos_current_mirror_0/IC Pmos_current_mirror_0/IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=2.2
X90 VDD Pmos_current_mirror_0/IA Pmos_current_mirror_0/IB VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=1 ps=6 w=1 l=2.2
X91 VDD VDD Pmos_current_mirror_0/IA VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=2.2
X92 VDD Pmos_current_mirror_0/IA Pmos_current_mirror_0/IC VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=2.2
X93 VDD Pmos_current_mirror_0/IA Pmos_current_mirror_0/IC VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=2.2
X94 VOUT Pmos_current_mirror_0/IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=2.2
X95 VOUT Pmos_current_mirror_0/IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=2.2
X96 VOUT Pmos_current_mirror_0/IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=2.2
X97 Pmos_current_mirror_0/IB Pmos_current_mirror_0/IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=2.2
X98 Pmos_current_mirror_0/IA Pmos_current_mirror_0/IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=2.2
X99 Pmos_current_mirror_0/IC Pmos_current_mirror_0/IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=2.2
X100 VDD Pmos_current_mirror_0/IA VOUT VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=2.2
X101 VDD Pmos_current_mirror_0/IA VOUT VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=2.2
X102 VDD Pmos_current_mirror_0/IA VOUT VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=2.2
X103 VDD Pmos_current_mirror_0/IA VOUT VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=2.2
X104 VDD Pmos_current_mirror_0/IA VOUT VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=2.2
X105 Pmos_current_mirror_0/IC Pmos_current_mirror_0/IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=2.2
X106 VDD VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=2.2
X107 Pmos_current_mirror_0/IC Pmos_current_mirror_0/IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=2.2
X108 VOUT Pmos_current_mirror_0/IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=2.2
X109 VOUT Pmos_current_mirror_0/IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=2.2
X110 VOUT Pmos_current_mirror_0/IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=2.2
X111 VOUT Pmos_current_mirror_0/IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=2.2
X112 VDD Pmos_current_mirror_0/IA VOUT VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=2.2
X113 VDD Pmos_current_mirror_0/IA VOUT VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=2.2
X114 VDD Pmos_current_mirror_0/IA Pmos_current_mirror_0/IC VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=2.2
X115 VDD Pmos_current_mirror_0/IA Pmos_current_mirror_0/IC VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=2.2
X116 m1_17410_n5244# Pmos_current_mirror_0/IB active_load_0/IA VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.35 pd=1.9 as=0.42 ps=3.4 w=1.4 l=2.6
X117 active_load_0/IA Pmos_current_mirror_0/IB m1_17410_n5244# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.4 as=0.35 ps=1.9 w=1.4 l=2.6
X118 Pmos_current_mirror_0/IA VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X119 Pmos_current_mirror_0/IB VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.3 ps=2.6 w=1 l=2
X120 VSS VSS Lower_Nmos_0/IA VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X121 VSS VSS Pmos_current_mirror_0/IB VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.3 pd=2.6 as=0.25 ps=1.5 w=1 l=2
X122 Pmos_current_mirror_0/IB Pmos_current_mirror_0/IB Lower_Nmos_0/IA VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X123 Lower_Nmos_0/IA VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X124 Lower_Nmos_0/IA Pmos_current_mirror_0/IB Pmos_current_mirror_0/IB VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X125 VSS VSS Pmos_current_mirror_0/IA VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X126 Pmos_current_mirror_0/IA Pmos_current_mirror_0/IB Lower_Nmos_0/IB VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X127 Lower_Nmos_0/IB Pmos_current_mirror_0/IB Pmos_current_mirror_0/IA VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X128 Pmos_current_mirror_0/IA VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=2 pd=12 as=0 ps=0 w=1 l=2
X129 Pmos_current_mirror_0/IB VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=2 pd=12 as=0 ps=0 w=1 l=2
X130 VSS VSS Lower_Nmos_0/IA VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=4 ps=24 w=1 l=2
X131 VSS VSS Pmos_current_mirror_0/IB VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=2
X132 Pmos_current_mirror_0/IB Pmos_current_mirror_0/IB Lower_Nmos_0/IA VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=2
X133 Lower_Nmos_0/IA VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=2
X134 Lower_Nmos_0/IA Pmos_current_mirror_0/IB Pmos_current_mirror_0/IB VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=2
X135 VSS VSS Pmos_current_mirror_0/IA VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=2
X136 Pmos_current_mirror_0/IA Pmos_current_mirror_0/IB Lower_Nmos_0/IB VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=6 ps=36 w=1 l=2
X137 Lower_Nmos_0/IB Pmos_current_mirror_0/IB Pmos_current_mirror_0/IA VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=2
X138 Lower_Nmos_0/IA Lower_Nmos_0/IA VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=3.2
X139 Lower_Nmos_0/IA VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.3 ps=2.6 w=1 l=3.2
X140 Lower_Nmos_0/IB VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=3.2
X141 VSS VSS Lower_Nmos_0/IA VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.3 pd=2.6 as=0.25 ps=1.5 w=1 l=3.2
X142 Lower_Nmos_0/IC Lower_Nmos_0/IA Lower_Nmos_0/IB VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=3.2
X143 Lower_Nmos_0/IC Lower_Nmos_0/IA Lower_Nmos_0/IB VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=3.2
X144 VSS Lower_Nmos_0/IA Lower_Nmos_0/IA VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=3.2
X145 Lower_Nmos_0/IB Lower_Nmos_0/IA Lower_Nmos_0/IC VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=3.2
X146 Lower_Nmos_0/IB Lower_Nmos_0/IA Lower_Nmos_0/IC VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=3.2
X147 Lower_Nmos_0/IC Lower_Nmos_0/IA Lower_Nmos_0/IB VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=3.2
X148 Lower_Nmos_0/IB Lower_Nmos_0/IA Lower_Nmos_0/IC VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=3.2
X149 Lower_Nmos_0/IB Lower_Nmos_0/IA Lower_Nmos_0/IC VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=3.2
X150 Lower_Nmos_0/IC Lower_Nmos_0/IA Lower_Nmos_0/IB VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=3.2
X151 VSS VSS Lower_Nmos_0/IB VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=3.2
X152 Lower_Nmos_0/IA Lower_Nmos_0/IA VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=3.2
X153 Lower_Nmos_0/IA VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.3 ps=2.6 w=1 l=3.2
X154 Lower_Nmos_0/IB VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=3.2
X155 VSS VSS Lower_Nmos_0/IA VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.3 pd=2.6 as=0.25 ps=1.5 w=1 l=3.2
X156 Lower_Nmos_0/IC Lower_Nmos_0/IA Lower_Nmos_0/IB VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=3.2
X157 Lower_Nmos_0/IC Lower_Nmos_0/IA Lower_Nmos_0/IB VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=3.2
X158 VSS Lower_Nmos_0/IA Lower_Nmos_0/IA VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=3.2
X159 Lower_Nmos_0/IB Lower_Nmos_0/IA Lower_Nmos_0/IC VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=3.2
X160 Lower_Nmos_0/IB Lower_Nmos_0/IA Lower_Nmos_0/IC VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=3.2
X161 Lower_Nmos_0/IC Lower_Nmos_0/IA Lower_Nmos_0/IB VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=3.2
X162 Lower_Nmos_0/IB Lower_Nmos_0/IA Lower_Nmos_0/IC VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=3.2
X163 Lower_Nmos_0/IB Lower_Nmos_0/IA Lower_Nmos_0/IC VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=3.2
X164 Lower_Nmos_0/IC Lower_Nmos_0/IA Lower_Nmos_0/IB VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=3.2
X165 VSS VSS Lower_Nmos_0/IB VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=3.2
X166 m1_17410_n5244# VOUT sky130_fd_pr__cap_mim_m3_1 l=8 w=8
X167 m1_17410_n5244# VOUT sky130_fd_pr__cap_mim_m3_1 l=8 w=8
X168 m1_17410_n5244# VOUT sky130_fd_pr__cap_mim_m3_1 l=8 w=8
X169 m1_17410_n5244# VOUT sky130_fd_pr__cap_mim_m3_1 l=8 w=8
C0 m1_17410_n5244# VOUT 29.48602f
C1 Pmos_current_mirror_0/IB VDD 2.21479f
C2 Pmos_current_mirror_0/IC Pmos_current_mirror_0/IA 3.2178f
C3 Lower_Nmos_0/IC Lower_Nmos_0/IA 4.67686f
C4 VOUT VDD 2.66933f
C5 Pmos_current_mirror_0/IC active_load_0/IA 3.7446f
C6 Pmos_current_mirror_0/IC VOUT 5.16991f
C7 active_load_0/IB Pmos_current_mirror_0/IC 3.62092f
C8 Vin+ Vin- 7.8812f
C9 Pmos_current_mirror_0/IB Pmos_current_mirror_0/IA 2.46011f
C10 Pmos_current_mirror_0/IC Vin- 4.1741f
C11 Pmos_current_mirror_0/IC VDD 2.33191f
C12 Lower_Nmos_0/IA Lower_Nmos_0/IB 6.14035f
C13 Pmos_current_mirror_0/IA VOUT 3.75574f
C14 Pmos_current_mirror_0/IC Vin+ 4.40894f
C15 VOUT active_load_0/IA 2.72808f
C16 active_load_0/IB active_load_0/IA 3.94623f
C17 Pmos_current_mirror_0/IA VDD 42.3693f
C18 m1_17410_n5244# VSS 4.27709f $ **FLOATING
C19 Lower_Nmos_0/IB VSS 3.18447f
C20 Lower_Nmos_0/IA VSS 33.08277f
C21 Lower_Nmos_0/IC VSS 3.21761f
C22 Pmos_current_mirror_0/IB VSS 17.06674f
C23 VOUT VSS 20.62634f
C24 Pmos_current_mirror_0/IA VSS 19.93994f
C25 VDD VSS 82.54808f
C26 Vin- VSS 2.91981f
C27 active_load_0/IA VSS 8.55239f
C28 Vin+ VSS 2.03204f
C29 Pmos_current_mirror_0/IC VSS 33.65339f
C30 active_load_0/IB VSS 11.94191f
.ends
