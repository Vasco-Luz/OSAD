* NGSPICE file created from Upper_Nmos.ext - technology: sky130A

.subckt Upper_Nmos VSS IF IA IB IE
X0 IA VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2 M=4
X1 IB VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.25 pd=1.5 as=0.3 ps=2.6 w=1 l=2 M=4
X2 VSS VSS IE VSS sky130_fd_pr__nfet_01v8_lvt ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2 M=4
X3 IB IB IE VSS sky130_fd_pr__nfet_01v8_lvt ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2 M=4
X4 IA IB IF VSS sky130_fd_pr__nfet_01v8_lvt ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2 M=4
C0 IB VSS 4.32532f
C1 IB 0 7.76271f
C2 VSS 0 7.75954f
.ends
