magic
tech sky130A
magscale 1 2
timestamp 1740487318
<< xpolycontact >>
rect -948 174 -878 606
rect -948 -606 -878 -174
rect -782 174 -712 606
rect -782 -606 -712 -174
rect -616 174 -546 606
rect -616 -606 -546 -174
rect -450 174 -380 606
rect -450 -606 -380 -174
rect -284 174 -214 606
rect -284 -606 -214 -174
rect -118 174 -48 606
rect -118 -606 -48 -174
rect 48 174 118 606
rect 48 -606 118 -174
rect 214 174 284 606
rect 214 -606 284 -174
rect 380 174 450 606
rect 380 -606 450 -174
rect 546 174 616 606
rect 546 -606 616 -174
rect 712 174 782 606
rect 712 -606 782 -174
rect 878 174 948 606
rect 878 -606 948 -174
<< ppolyres >>
rect -948 -174 -878 174
rect -782 -174 -712 174
rect -616 -174 -546 174
rect -450 -174 -380 174
rect -284 -174 -214 174
rect -118 -174 -48 174
rect 48 -174 118 174
rect 214 -174 284 174
rect 380 -174 450 174
rect 546 -174 616 174
rect 712 -174 782 174
rect 878 -174 948 174
<< viali >>
rect -932 191 -894 588
rect -766 191 -728 588
rect -600 191 -562 588
rect -434 191 -396 588
rect -268 191 -230 588
rect -102 191 -64 588
rect 64 191 102 588
rect 230 191 268 588
rect 396 191 434 588
rect 562 191 600 588
rect 728 191 766 588
rect 894 191 932 588
rect -932 -588 -894 -191
rect -766 -588 -728 -191
rect -600 -588 -562 -191
rect -434 -588 -396 -191
rect -268 -588 -230 -191
rect -102 -588 -64 -191
rect 64 -588 102 -191
rect 230 -588 268 -191
rect 396 -588 434 -191
rect 562 -588 600 -191
rect 728 -588 766 -191
rect 894 -588 932 -191
<< metal1 >>
rect -938 588 -888 600
rect -938 191 -932 588
rect -894 191 -888 588
rect -938 179 -888 191
rect -772 588 -722 600
rect -772 191 -766 588
rect -728 191 -722 588
rect -772 179 -722 191
rect -606 588 -556 600
rect -606 191 -600 588
rect -562 191 -556 588
rect -606 179 -556 191
rect -440 588 -390 600
rect -440 191 -434 588
rect -396 191 -390 588
rect -440 179 -390 191
rect -274 588 -224 600
rect -274 191 -268 588
rect -230 191 -224 588
rect -274 179 -224 191
rect -108 588 -58 600
rect -108 191 -102 588
rect -64 191 -58 588
rect -108 179 -58 191
rect 58 588 108 600
rect 58 191 64 588
rect 102 191 108 588
rect 58 179 108 191
rect 224 588 274 600
rect 224 191 230 588
rect 268 191 274 588
rect 224 179 274 191
rect 390 588 440 600
rect 390 191 396 588
rect 434 191 440 588
rect 390 179 440 191
rect 556 588 606 600
rect 556 191 562 588
rect 600 191 606 588
rect 556 179 606 191
rect 722 588 772 600
rect 722 191 728 588
rect 766 191 772 588
rect 722 179 772 191
rect 888 588 938 600
rect 888 191 894 588
rect 932 191 938 588
rect 888 179 938 191
rect -938 -191 -888 -179
rect -938 -588 -932 -191
rect -894 -588 -888 -191
rect -938 -600 -888 -588
rect -772 -191 -722 -179
rect -772 -588 -766 -191
rect -728 -588 -722 -191
rect -772 -600 -722 -588
rect -606 -191 -556 -179
rect -606 -588 -600 -191
rect -562 -588 -556 -191
rect -606 -600 -556 -588
rect -440 -191 -390 -179
rect -440 -588 -434 -191
rect -396 -588 -390 -191
rect -440 -600 -390 -588
rect -274 -191 -224 -179
rect -274 -588 -268 -191
rect -230 -588 -224 -191
rect -274 -600 -224 -588
rect -108 -191 -58 -179
rect -108 -588 -102 -191
rect -64 -588 -58 -191
rect -108 -600 -58 -588
rect 58 -191 108 -179
rect 58 -588 64 -191
rect 102 -588 108 -191
rect 58 -600 108 -588
rect 224 -191 274 -179
rect 224 -588 230 -191
rect 268 -588 274 -191
rect 224 -600 274 -588
rect 390 -191 440 -179
rect 390 -588 396 -191
rect 434 -588 440 -191
rect 390 -600 440 -588
rect 556 -191 606 -179
rect 556 -588 562 -191
rect 600 -588 606 -191
rect 556 -600 606 -588
rect 722 -191 772 -179
rect 722 -588 728 -191
rect 766 -588 772 -191
rect 722 -600 772 -588
rect 888 -191 938 -179
rect 888 -588 894 -191
rect 932 -588 938 -191
rect 888 -600 938 -588
<< properties >>
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 1.9 m 1 nx 12 wmin 0.350 lmin 0.50 class resistor rho 319.8 val 2.849k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
