magic
tech sky130A
magscale 1 2
timestamp 1693703138
<< locali >>
rect 116 126 152 1118
rect 188 976 298 1120
rect 2586 978 2696 1122
rect 2732 126 2768 1134
rect 74 -476 108 -226
rect 152 -376 248 -232
rect 2550 -376 2646 -232
rect 2690 -446 2724 -222
<< viali >>
rect 1292 1102 1590 1142
rect 1210 -2156 1582 -2120
<< metal1 >>
rect 1410 1160 1470 1280
rect 1282 1142 1602 1160
rect 1282 1102 1292 1142
rect 1590 1102 1602 1142
rect 1282 1100 1602 1102
rect 328 1064 2556 1100
rect 328 898 376 1064
rect 420 1030 502 1036
rect 420 978 426 1030
rect 496 978 502 1030
rect 420 972 502 978
rect 638 1030 720 1036
rect 638 978 644 1030
rect 714 978 720 1030
rect 638 972 720 978
rect 764 904 812 1064
rect 856 1030 938 1036
rect 856 978 862 1030
rect 932 978 938 1030
rect 856 972 938 978
rect 1074 1030 1156 1036
rect 1074 978 1080 1030
rect 1150 978 1156 1030
rect 1074 972 1156 978
rect 1200 904 1248 1064
rect 1292 1030 1374 1036
rect 1292 978 1298 1030
rect 1368 978 1374 1030
rect 1292 972 1374 978
rect 1510 1030 1592 1036
rect 1510 978 1516 1030
rect 1586 978 1592 1030
rect 1510 972 1592 978
rect 1636 904 1684 1064
rect 1728 1030 1810 1036
rect 1728 978 1734 1030
rect 1804 978 1810 1030
rect 1728 972 1810 978
rect 1946 1030 2028 1036
rect 1946 978 1952 1030
rect 2022 978 2028 1030
rect 1946 972 2028 978
rect 2072 910 2120 1064
rect 2164 1030 2246 1036
rect 2164 978 2170 1030
rect 2240 978 2246 1030
rect 2164 972 2246 978
rect 2382 1030 2464 1036
rect 2382 978 2388 1030
rect 2458 978 2464 1030
rect 2382 972 2464 978
rect 2508 900 2556 1064
rect 546 70 594 172
rect 982 70 1030 178
rect 1418 70 1466 178
rect 1854 70 1902 174
rect 2290 70 2338 176
rect 546 32 2338 70
rect 1376 -260 1422 32
rect 1854 30 1902 32
rect 286 -290 2512 -260
rect 286 -440 332 -290
rect 380 -324 456 -318
rect 380 -376 386 -324
rect 450 -376 456 -324
rect 380 -382 456 -376
rect 598 -324 674 -318
rect 598 -376 604 -324
rect 668 -376 674 -324
rect 598 -382 674 -376
rect 722 -416 768 -290
rect 816 -324 892 -318
rect 816 -376 822 -324
rect 886 -376 892 -324
rect 816 -382 892 -376
rect 1034 -324 1110 -318
rect 1034 -376 1040 -324
rect 1104 -376 1110 -324
rect 1034 -382 1110 -376
rect 1158 -420 1204 -290
rect 1252 -324 1328 -318
rect 1252 -376 1258 -324
rect 1322 -376 1328 -324
rect 1252 -382 1328 -376
rect 1470 -324 1546 -318
rect 1470 -376 1476 -324
rect 1540 -376 1546 -324
rect 1470 -382 1546 -376
rect 1594 -420 1640 -290
rect 1688 -324 1764 -318
rect 1688 -376 1694 -324
rect 1758 -376 1764 -324
rect 1688 -382 1764 -376
rect 1906 -324 1982 -318
rect 1906 -376 1912 -324
rect 1976 -376 1982 -324
rect 1906 -382 1982 -376
rect 2030 -424 2076 -290
rect 2124 -324 2200 -318
rect 2124 -376 2130 -324
rect 2194 -376 2200 -324
rect 2124 -382 2200 -376
rect 2342 -324 2418 -318
rect 2342 -376 2348 -324
rect 2412 -376 2418 -324
rect 2342 -382 2418 -376
rect 2466 -432 2512 -290
rect 504 -2080 550 -1970
rect 940 -2080 986 -1990
rect 1376 -2080 1422 -1992
rect 1812 -2080 1858 -1990
rect 2248 -2080 2294 -1992
rect 504 -2110 2294 -2080
rect 1158 -2120 1640 -2110
rect 1158 -2156 1210 -2120
rect 1582 -2156 1640 -2120
rect 1158 -2162 1640 -2156
rect 1322 -2258 1464 -2162
<< via1 >>
rect 426 978 496 1030
rect 644 978 714 1030
rect 862 978 932 1030
rect 1080 978 1150 1030
rect 1298 978 1368 1030
rect 1516 978 1586 1030
rect 1734 978 1804 1030
rect 1952 978 2022 1030
rect 2170 978 2240 1030
rect 2388 978 2458 1030
rect 386 -376 450 -324
rect 604 -376 668 -324
rect 822 -376 886 -324
rect 1040 -376 1104 -324
rect 1258 -376 1322 -324
rect 1476 -376 1540 -324
rect 1694 -376 1758 -324
rect 1912 -376 1976 -324
rect 2130 -376 2194 -324
rect 2348 -376 2412 -324
<< metal2 >>
rect -136 1036 1342 1038
rect -136 1030 2464 1036
rect -136 978 426 1030
rect 496 978 644 1030
rect 714 978 862 1030
rect 932 978 1080 1030
rect 1150 978 1298 1030
rect 1368 978 1516 1030
rect 1586 978 1734 1030
rect 1804 978 1952 1030
rect 2022 978 2170 1030
rect 2240 978 2388 1030
rect 2458 978 2464 1030
rect -136 972 2464 978
rect -136 970 1342 972
rect -134 -324 2418 -318
rect -134 -376 386 -324
rect 450 -376 604 -324
rect 668 -376 822 -324
rect 886 -376 1040 -324
rect 1104 -376 1258 -324
rect 1322 -376 1476 -324
rect 1540 -376 1694 -324
rect 1758 -376 1912 -324
rect 1976 -376 2130 -324
rect 2194 -376 2348 -324
rect 2412 -376 2418 -324
rect -134 -382 2418 -376
use sky130_fd_pr__nfet_g5v0d10v5_4HWKKE  sky130_fd_pr__nfet_g5v0d10v5_4HWKKE_0
timestamp 1693700175
transform 1 0 1399 0 1 -1183
box -1507 -1027 1507 1027
use sky130_fd_pr__pfet_g5v0d10v5_CHJVJW  sky130_fd_pr__pfet_g5v0d10v5_CHJVJW_0
timestamp 1693699723
transform 1 0 1442 0 1 567
box -1537 -662 1537 662
<< labels >>
flabel metal1 1410 1142 1470 1280 0 FreeSans 1600 0 0 0 VDD
port 1 nsew
flabel metal1 1322 -2258 1464 -2156 0 FreeSans 1600 0 0 0 VSS
port 3 nsew
flabel metal2 -134 -382 386 -318 0 FreeSans 1600 0 0 0 VIN
port 5 nsew
flabel metal1 1376 -290 1422 70 0 FreeSans 1600 0 0 0 VOUT
port 7 nsew
flabel metal2 -136 970 426 1038 0 FreeSans 1600 0 0 0 VB
port 9 nsew
<< end >>
