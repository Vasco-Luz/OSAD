** sch_path: /home/gim/Desktop/OSAD/my_ip/testbenches_sky/single_ended_OTAS_testbenches/single_ended_OTA_AC_TB.sch
**.subckt single_ended_OTA_AC_TB
*  x1 -  UUT  IS MISSING !!!!
V1 VDD GND VDD
V2 VSS GND VSS
V4 VIN+ net1 ac 0.5
V6 net2 net1 V_OFF
V3 net1 GND VCM
V5 VIN- net2 ac -0.5
C1 VOUT VSS CL m=1
*  x2 -  UUT  IS MISSING !!!!
C2 VOUT_cm VSS CL m=1
V8 net4 net3 V_OFF
V9 net10 GND VCM
V7 net3 net10 ac 1
*  x3 -  UUT  IS MISSING !!!!
C3 VOUT_a- VSS CL m=1
V10 net6 net5 V_OFF
V11 net5 GND VCM
V13 net7 VSS ac 1
*  x4 -  UUT  IS MISSING !!!!
C4 VOUT_a+ VSS CL m=1
V12 net9 net8 V_OFF
V14 net8 GND VCM
V15 net11 VDD ac 1
**** begin user architecture code
.lib /home/gim/PDK/sky130A/libs.tech/combined/sky130.lib.spice tt


.Temp 27
.param VDD = 1.8
.param VSS = 0
.param VCM={(VDD-VSS)/2}
.param VCM_NEG={-VCM}
.param V_OFF = 12.93u
.param CL = 3p

.control
save all

ac dec 100 1 10G
wrdata VIN_sweep_AC.csv db(v(VOUT)) phase(VOUT) db(v(VOUT_cm)) db(v(VOUT_a-)) db(v(VOUT_a+))
plot db(v(VOUT)) phase(VOUT)
plot db(v(VOUT_cm))
plot db(v(VOUT_a-))
plot db(v(VOUT_a+))

.endc

**** end user architecture code
**.ends
.GLOBAL GND
.end
