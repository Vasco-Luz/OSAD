** sch_path: /foss/designs/OSAD/Learning/single_ended_amplifiers/Design_and_Analysis_of_Two-Stage_CMOS_Operational_Amplifier_for_Fluorescence_Signal_Processing_sky130_5V/amplifier_design/OTA_DC_TB.sch
**.subckt OTA_DC_TB
V1 VDD GND VDD
V2 VSS GND VSS
V4 VIN+ VSS 2.5
Vmeas VDD net1 0
.save i(vmeas)
x1 net1 VSS VOUT VIN+ VOUT UUT_VA_sky
**** begin user architecture code
.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice tt

.Temp 27
.param VDD = 5
.param VSS = 0

.control
save all
dc V4 0 5 0.01
wrdata VIN_sweep_DC.csv v(VOUT) i(Vmeas)
plot v(VOUT) v(VIN+)
plot i(Vmeas)

.endc

**** end user architecture code
**.ends

* expanding   symbol:  Sky130A/UUT_sky/UUT_VA_sky.sym # of pins=5
** sym_path: /foss/designs/OSAD/my_ip/LIB/Sky130A/UUT_sky/UUT_VA_sky.sym
** sch_path: /foss/designs/OSAD/my_ip/LIB/Sky130A/UUT_sky/UUT_VA_sky.sch
.subckt UUT_VA_sky VDD VSS VIN- VIN+ VOUT
*.iopin VDD
*.iopin VSS
*.iopin VIN-
*.iopin VIN+
*.iopin VOUT
x1 VDD VSS VIN+ VIN- VOUT A001
.ends


* expanding   symbol:
*+  Sky130A/Learning/Design_of_Two-Stage_CMOS_Operational_Amplifier_for_Fluorescence_Signal_Processing_5V/A001.sym # of pins=5
** sym_path: /foss/designs/OSAD/my_ip/LIB/Sky130A/Learning/Design_of_Two-Stage_CMOS_Operational_Amplifier_for_Fluorescence_Signal_Processing_5V/A001.sym
** sch_path: /foss/designs/OSAD/my_ip/LIB/Sky130A/Learning/Design_of_Two-Stage_CMOS_Operational_Amplifier_for_Fluorescence_Signal_Processing_5V/A001.sch
.subckt A001 VDD VSS Vin+ Vin- VOUT
*.iopin VDD
*.iopin VSS
*.iopin Vin+
*.iopin Vin-
*.iopin VOUT
XM5 VB2 VB1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2.2 W='1 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=2
+ m=2
XM6 VB1 VB1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2.2 W='1 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=2
+ m=2
XR2 VSS net2 VSS sky130_fd_pr__res_high_po_0p35 L=20.4 mult=1 m=1
XM7 net1 net1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=3.2 W='1 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=2
+ m=2
XM8 net3 net1 net2 VSS sky130_fd_pr__nfet_g5v0d10v5 L=3.2 W='1 * 8 ' nf=8 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=2
+ m=2
XM9 VB1 VB2 net3 VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W='1 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=2
+ m=2
XM10 VB2 VB2 net1 VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W='1 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=2
+ m=2
XM1 net4 VB1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2.2 W='1 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=8
+ m=8
XM2 VOUT VB1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2.2 W='1 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=16
+ m=16
XM3 net6 Vin- net4 net4 sky130_fd_pr__pfet_g5v0d10v5 L=1 W='4 * 4 ' nf=4 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=4
+ m=4
XM4 net5 Vin+ net4 net4 sky130_fd_pr__pfet_g5v0d10v5 L=1 W='4 * 4 ' nf=4 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=4
+ m=4
XM11 net5 net6 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W='1 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=2
+ m=2
XM12 net6 net6 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W='1 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=2
+ m=2
XM13 VOUT net5 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W='4 * 4 ' nf=4 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=2
+ m=2
XM14 net7 VB2 net5 VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W='1 * 1 ' nf=1 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=2
+ m=2
XC1 VOUT net7 sky130_fd_pr__cap_mim_m3_1 W=8 L=8 MF=4 m=4
.ends

.GLOBAL GND
.end
