magic
tech sky130A
magscale 1 2
timestamp 1738951789
<< nwell >>
rect -753 -216 793 236
rect -723 -244 793 -216
rect -723 -250 723 -244
<< mvpmos >>
rect -629 -150 -29 150
rect 29 -150 629 150
<< mvpdiff >>
rect -687 138 -629 150
rect -687 -138 -675 138
rect -641 -138 -629 138
rect -687 -150 -629 -138
rect -29 138 29 150
rect -29 -138 -17 138
rect 17 -138 29 138
rect -29 -150 29 -138
rect 629 138 687 150
rect 629 -138 641 138
rect 675 -138 687 138
rect 629 -150 687 -138
<< mvpdiffc >>
rect -675 -138 -641 138
rect -17 -138 17 138
rect 641 -138 675 138
<< poly >>
rect -629 150 -29 186
rect 29 150 629 186
rect -629 -197 -29 -150
rect -629 -214 -556 -197
rect -572 -231 -556 -214
rect -102 -214 -29 -197
rect 29 -197 629 -150
rect 29 -214 102 -197
rect -102 -231 -86 -214
rect -572 -247 -86 -231
rect 86 -231 102 -214
rect 556 -214 629 -197
rect 556 -231 572 -214
rect 86 -247 572 -231
<< polycont >>
rect -556 -231 -102 -197
rect 102 -231 556 -197
<< locali >>
rect -675 138 -641 154
rect -675 -154 -641 -138
rect -17 138 17 154
rect -17 -154 17 -138
rect 641 138 675 154
rect 641 -154 675 -138
rect -572 -231 -556 -197
rect -102 -231 -86 -197
rect 86 -231 102 -197
rect 556 -231 572 -197
<< viali >>
rect -675 -138 -641 138
rect -17 -138 17 138
rect 641 -138 675 138
rect -556 -231 -102 -197
rect 102 -231 556 -197
<< metal1 >>
rect -681 138 -635 150
rect -681 -138 -675 138
rect -641 -138 -635 138
rect -681 -150 -635 -138
rect -23 138 23 150
rect -23 -138 -17 138
rect 17 -138 23 138
rect -23 -150 23 -138
rect 635 138 681 150
rect 635 -138 641 138
rect 675 -138 681 138
rect 635 -150 681 -138
rect -568 -197 -90 -191
rect -568 -231 -556 -197
rect -102 -231 -90 -197
rect -568 -237 -90 -231
rect 90 -197 568 -191
rect 90 -231 102 -197
rect 556 -231 568 -197
rect 90 -237 568 -231
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1.5 l 3 m 1 nf 2 diffcov 100 polycov 80 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 1 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 80 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
