** sch_path: /foss/designs/OSAD/Learning/single_ended_amplifiers/Design_and_Analysis_of_Two-Stage_CMOS_Operational_Amplifier_for_Fluorescence_Signal_Processing_sky130_5V/transimpedance_cell_design/transcondutance_cell_design.sch
**.subckt transcondutance_cell_design
V1 VDD GND VDD
V2 VSS GND VSS
XR6 VSS net11 VSS sky130_fd_pr__res_high_po_0p35 L=30 mult=1 m=1
R1 net3 net2 0.001 m=1
G1 net5 net1 net3 net2 1000
Vmeas net4 net3 0
.save i(vmeas)
Vmeas1 net4 net5 0
.save i(vmeas1)
V3 net4 GND 1.8
XM1 net2 net1 net11 VSS sky130_fd_pr__nfet_g5v0d10v5 L=4 W='0.6 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=8
+ m=8
XM2 net1 net1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=4 W='0.6 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=2
+ m=2
G2 net6 VSS net3 net2 1000
XM4 net6 net6 net4 net4 sky130_fd_pr__pfet_g5v0d10v5 L=3 W='1.5 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=2
+ m=2
XM3 net7 net6 net4 net4 sky130_fd_pr__pfet_g5v0d10v5 L=3 W='1.5 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=2
+ m=2
Vmeas2 net7 VSS 0
.save i(vmeas2)
XM5 net8 net8 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=3 W='1.5 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=2
+ m=2
XM6 net15 net8 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=3 W='1.5 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=2
+ m=2
XM7 net12 net9 net10 VSS sky130_fd_pr__nfet_g5v0d10v5 L=4 W='0.6 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=8
+ m=8
XM8 net9 net9 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=4 W='0.6 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=2
+ m=2
XM9 net14 net13 net12 VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W='0.6 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=2
+ m=2
XM10 net13 net13 net9 VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W='0.6 * 2 ' nf=2 ad='int((nf+1)/2) * W / nf * 0.29' as='int((nf+2)/2) * W / nf * 0.29'
+ pd='2*int((nf+1)/2) * (W / nf + 0.29)' ps='2*int((nf+2)/2) * (W / nf + 0.29)' nrd='0.29 / W ' nrs='0.29 / W ' sa=0 sb=0 sd=0 mult=2
+ m=2
Vmeas3 net8 net14 0
.save i(vmeas3)
Vmeas4 net15 net13 0
.save i(vmeas4)
XR2 VSS net10 VSS sky130_fd_pr__res_high_po_0p35 L=30 mult=1 m=1
**** begin user architecture code
.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice tt_mm


.Temp 27
.param VDD = 5
.param VSS = 0


.control
save all

save

dc Temp -40 125 1
plot i(Vmeas1) i(Vmeas2)
plot i(Vmeas3) i(Vmeas4)
wrdata data.csv i(Vmeas3) i(Vmeas4)


op
print i(Vmeas1)
print v(net2)




.endc

**** end user architecture code
**.ends
.GLOBAL GND
.end
