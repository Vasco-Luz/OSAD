magic
tech sky130A
magscale 1 2
timestamp 1738972435
<< nwell >>
rect -887 -447 887 447
<< mvpmos >>
rect -629 -150 -29 150
rect 29 -150 629 150
<< mvpdiff >>
rect -687 138 -629 150
rect -687 -138 -675 138
rect -641 -138 -629 138
rect -687 -150 -629 -138
rect -29 138 29 150
rect -29 -138 -17 138
rect 17 -138 29 138
rect -29 -150 29 -138
rect 629 138 687 150
rect 629 -138 641 138
rect 675 -138 687 138
rect 629 -150 687 -138
<< mvpdiffc >>
rect -675 -138 -641 138
rect -17 -138 17 138
rect 641 -138 675 138
<< mvnsubdiff >>
rect -821 369 821 381
rect -821 335 -713 369
rect 713 335 821 369
rect -821 323 821 335
rect -821 273 -763 323
rect -821 -273 -809 273
rect -775 -273 -763 273
rect 763 273 821 323
rect -821 -323 -763 -273
rect 763 -273 775 273
rect 809 -273 821 273
rect 763 -323 821 -273
rect -821 -335 821 -323
rect -821 -369 -713 -335
rect 713 -369 821 -335
rect -821 -381 821 -369
<< mvnsubdiffcont >>
rect -713 335 713 369
rect -809 -273 -775 273
rect 775 -273 809 273
rect -713 -369 713 -335
<< poly >>
rect -629 231 -29 247
rect -629 197 -613 231
rect -45 197 -29 231
rect -629 150 -29 197
rect 29 231 629 247
rect 29 197 45 231
rect 613 197 629 231
rect 29 150 629 197
rect -629 -197 -29 -150
rect -629 -231 -613 -197
rect -45 -231 -29 -197
rect -629 -247 -29 -231
rect 29 -197 629 -150
rect 29 -231 45 -197
rect 613 -231 629 -197
rect 29 -247 629 -231
<< polycont >>
rect -613 197 -45 231
rect 45 197 613 231
rect -613 -231 -45 -197
rect 45 -231 613 -197
<< locali >>
rect -809 335 -713 369
rect 713 335 809 369
rect -809 273 -775 335
rect 775 273 809 335
rect -629 197 -613 231
rect -45 197 -29 231
rect 29 197 45 231
rect 613 197 629 231
rect -675 138 -641 154
rect -675 -154 -641 -138
rect -17 138 17 154
rect -17 -154 17 -138
rect 641 138 675 154
rect 641 -154 675 -138
rect -629 -231 -613 -197
rect -45 -231 -29 -197
rect 29 -231 45 -197
rect 613 -231 629 -197
rect -809 -335 -775 -273
rect 775 -335 809 -273
rect -809 -369 -713 -335
rect 713 -369 809 -335
<< viali >>
rect -613 197 -45 231
rect 45 197 613 231
rect -675 -138 -641 138
rect -17 -138 17 138
rect 641 -138 675 138
rect -613 -231 -45 -197
rect 45 -231 613 -197
<< metal1 >>
rect -625 231 -33 237
rect -625 197 -613 231
rect -45 197 -33 231
rect -625 191 -33 197
rect 33 231 625 237
rect 33 197 45 231
rect 613 197 625 231
rect 33 191 625 197
rect -681 138 -635 150
rect -681 -138 -675 138
rect -641 -138 -635 138
rect -681 -150 -635 -138
rect -23 138 23 150
rect -23 -138 -17 138
rect 17 -138 23 138
rect -23 -150 23 -138
rect 635 138 681 150
rect 635 -138 641 138
rect 675 -138 681 138
rect 635 -150 681 -138
rect -625 -197 -33 -191
rect -625 -231 -613 -197
rect -45 -231 -33 -197
rect -625 -237 -33 -231
rect 33 -197 625 -191
rect 33 -231 45 -197
rect 613 -231 625 -197
rect 33 -237 625 -231
<< properties >>
string FIXED_BBOX -792 -352 792 352
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1.5 l 3 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
