magic
tech sky130a
timestamp 1739287221
<< checkpaint >>
rect -47 -88 407 204
<< l65d20 >>
rect 0 0 360 150
<< l66d44 >>
rect 337 13 354 30
rect 337 49 354 66
rect 337 85 354 102
rect 337 121 354 138
rect 46 -45 63 -28
rect 82 -45 99 -28
rect 118 -45 135 -28
rect 154 -45 171 -28
rect 190 -45 207 -28
rect 226 -45 243 -28
rect 262 -45 279 -28
rect 298 -45 315 -28
rect 7 13 24 30
rect 7 49 24 66
rect 7 85 24 102
rect 7 121 24 138
<< l67d20 >>
rect 337 5 354 146
rect 38 -45 323 -28
rect 7 5 24 146
<< l67d44 >>
rect 337 13 354 30
rect 337 49 354 66
rect 337 85 354 102
rect 337 121 354 138
rect 46 -45 63 -28
rect 82 -45 99 -28
rect 118 -45 135 -28
rect 154 -45 171 -28
rect 190 -45 207 -28
rect 226 -45 243 -28
rect 262 -45 279 -28
rect 298 -45 315 -28
rect 7 13 24 30
rect 7 49 24 66
rect 7 85 24 102
rect 7 121 24 138
<< l68d20 >>
rect 334 7 357 144
rect 40 -48 321 -25
rect 4 7 27 144
<< l66d20 >>
rect 30 -53 330 -20
rect 30 -20 330 170
<< l95d20 >>
rect 29 -54 331 -19
<< l94d20 >>
rect -13 -13 373 163
<< l64d20 >>
rect -47 -88 407 204
<< l75d20 >>
rect -47 -88 407 204
<< end >>
