** sch_path: /foss/designs/OSAD/Learning/fully_differencial/Indirect_Compensation_Techniques_for_Three_Stage_Fully_Differential_Op_amps_IHP130/testbenches/transimpedance_cell_tb_.sch
**.subckt transimpedance_cell_tb_
XR1 net1 VDD rhigh w=0.5e-6 l=5.85e-6 m=1 b=0
R2 net2 VSS 0.001 m=1
G1 net3 net4 net2 VSS 1000
V1 VDD GND VDD
V2 VSS GND VSS
XM1 net2 net3 net1 VDD sg13_hv_pmos w=2.0u l=3u ng=2 m=8
XM2 net3 net3 VDD VDD sg13_hv_pmos w=2.0u l=3u ng=2 m=2
Vmeas net4 VSS 0
.save i(vmeas)
G2 VDD net5 net2 VSS 1000
XM3 net5 net5 VSS VSS sg13_hv_nmos w=4.5u l=2u ng=2 m=2
Vmeas1 net7 net6 0
.save i(vmeas1)
V3 net7 GND 1.65
XM4 net6 net5 VSS VSS sg13_hv_nmos w=4.5u l=2u ng=2 m=2
XM6 net8 net9 VSS VSS sg13_hv_nmos w=4.5u l=2u ng=2 m=2
Vmeas2 VDD net8 0
.save i(vmeas2)
x1 VDD VSS net9 bias_cell
**** begin user architecture code


.param mm_ok=1
.param mc_ok=1
.param temp=27
.param VDD=3.3
.param VSS=0
.control
	save all
	dc V3 0 3.3 0.01
	plot i(Vmeas1)
	op
	dc temp -40 125 1
	plot i(Vmeas2)
	write op.raw
.endc



.lib cornerMOShv.lib mos_tt


.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerRES.lib res_typ

**** end user architecture code
**.ends

* expanding   symbol:  ihp-sg13g2/FD_opamp001/bias_cell.sym # of pins=3
** sym_path: /foss/designs/OSAD/my_ip/LIB/ihp-sg13g2/FD_opamp001/bias_cell.sym
** sch_path: /foss/designs/OSAD/my_ip/LIB/ihp-sg13g2/FD_opamp001/bias_cell.sch
.subckt bias_cell VDD VSS VB
*.iopin VDD
*.iopin VSS
*.iopin VB
XM5 net4 VB VSS VSS sg13_hv_nmos w=4.5u l=2u ng=2 m=2
XM6 VB VB VSS VSS sg13_hv_nmos w=4.5u l=2u ng=2 m=2
XR3 net1 VDD rhigh w=0.5e-6 l=1.95e-6 m=1 b=0
XM7 net3 net2 net1 VDD sg13_hv_pmos w=2.0u l=3u ng=2 m=8
XM8 net2 net2 VDD VDD sg13_hv_pmos w=2.0u l=3u ng=2 m=2
XM9 net4 net4 net2 VDD sg13_hv_pmos w=2.0u l=3u ng=2 m=2
XM10 net5 net4 net3 VDD sg13_hv_pmos w=2.0u l=3u ng=2 m=2
Vmeas2 net5 VB 0
.save i(vmeas2)
.ends

.GLOBAL GND
.end
