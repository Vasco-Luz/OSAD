magic
tech sky130A
magscale 1 2
timestamp 1693700175
<< pwell >>
rect -1507 -1058 1507 1058
<< mvnmos >>
rect -1279 -800 -1119 800
rect -1061 -800 -901 800
rect -843 -800 -683 800
rect -625 -800 -465 800
rect -407 -800 -247 800
rect -189 -800 -29 800
rect 29 -800 189 800
rect 247 -800 407 800
rect 465 -800 625 800
rect 683 -800 843 800
rect 901 -800 1061 800
rect 1119 -800 1279 800
<< mvndiff >>
rect -1337 788 -1279 800
rect -1337 -788 -1325 788
rect -1291 -788 -1279 788
rect -1337 -800 -1279 -788
rect -1119 788 -1061 800
rect -1119 -788 -1107 788
rect -1073 -788 -1061 788
rect -1119 -800 -1061 -788
rect -901 788 -843 800
rect -901 -788 -889 788
rect -855 -788 -843 788
rect -901 -800 -843 -788
rect -683 788 -625 800
rect -683 -788 -671 788
rect -637 -788 -625 788
rect -683 -800 -625 -788
rect -465 788 -407 800
rect -465 -788 -453 788
rect -419 -788 -407 788
rect -465 -800 -407 -788
rect -247 788 -189 800
rect -247 -788 -235 788
rect -201 -788 -189 788
rect -247 -800 -189 -788
rect -29 788 29 800
rect -29 -788 -17 788
rect 17 -788 29 788
rect -29 -800 29 -788
rect 189 788 247 800
rect 189 -788 201 788
rect 235 -788 247 788
rect 189 -800 247 -788
rect 407 788 465 800
rect 407 -788 419 788
rect 453 -788 465 788
rect 407 -800 465 -788
rect 625 788 683 800
rect 625 -788 637 788
rect 671 -788 683 788
rect 625 -800 683 -788
rect 843 788 901 800
rect 843 -788 855 788
rect 889 -788 901 788
rect 843 -800 901 -788
rect 1061 788 1119 800
rect 1061 -788 1073 788
rect 1107 -788 1119 788
rect 1061 -800 1119 -788
rect 1279 788 1337 800
rect 1279 -788 1291 788
rect 1325 -788 1337 788
rect 1279 -800 1337 -788
<< mvndiffc >>
rect -1325 -788 -1291 788
rect -1107 -788 -1073 788
rect -889 -788 -855 788
rect -671 -788 -637 788
rect -453 -788 -419 788
rect -235 -788 -201 788
rect -17 -788 17 788
rect 201 -788 235 788
rect 419 -788 453 788
rect 637 -788 671 788
rect 855 -788 889 788
rect 1073 -788 1107 788
rect 1291 -788 1325 788
<< mvpsubdiff >>
rect -1471 1010 1471 1022
rect -1471 976 -1363 1010
rect 1363 976 1471 1010
rect -1471 964 1471 976
rect -1471 914 -1413 964
rect -1471 -914 -1459 914
rect -1425 -914 -1413 914
rect 1413 914 1471 964
rect -1471 -964 -1413 -914
rect 1413 -914 1425 914
rect 1459 -914 1471 914
rect 1413 -964 1471 -914
rect -1471 -976 1471 -964
rect -1471 -1010 -1363 -976
rect 1363 -1010 1471 -976
rect -1471 -1022 1471 -1010
<< mvpsubdiffcont >>
rect -1363 976 1363 1010
rect -1459 -914 -1425 914
rect 1425 -914 1459 914
rect -1363 -1010 1363 -976
<< poly >>
rect -1279 872 -1119 888
rect -1279 838 -1263 872
rect -1135 838 -1119 872
rect -1279 800 -1119 838
rect -1061 872 -901 888
rect -1061 838 -1045 872
rect -917 838 -901 872
rect -1061 800 -901 838
rect -843 872 -683 888
rect -843 838 -827 872
rect -699 838 -683 872
rect -843 800 -683 838
rect -625 872 -465 888
rect -625 838 -609 872
rect -481 838 -465 872
rect -625 800 -465 838
rect -407 872 -247 888
rect -407 838 -391 872
rect -263 838 -247 872
rect -407 800 -247 838
rect -189 872 -29 888
rect -189 838 -173 872
rect -45 838 -29 872
rect -189 800 -29 838
rect 29 872 189 888
rect 29 838 45 872
rect 173 838 189 872
rect 29 800 189 838
rect 247 872 407 888
rect 247 838 263 872
rect 391 838 407 872
rect 247 800 407 838
rect 465 872 625 888
rect 465 838 481 872
rect 609 838 625 872
rect 465 800 625 838
rect 683 872 843 888
rect 683 838 699 872
rect 827 838 843 872
rect 683 800 843 838
rect 901 872 1061 888
rect 901 838 917 872
rect 1045 838 1061 872
rect 901 800 1061 838
rect 1119 872 1279 888
rect 1119 838 1135 872
rect 1263 838 1279 872
rect 1119 800 1279 838
rect -1279 -838 -1119 -800
rect -1279 -872 -1263 -838
rect -1135 -872 -1119 -838
rect -1279 -888 -1119 -872
rect -1061 -838 -901 -800
rect -1061 -872 -1045 -838
rect -917 -872 -901 -838
rect -1061 -888 -901 -872
rect -843 -838 -683 -800
rect -843 -872 -827 -838
rect -699 -872 -683 -838
rect -843 -888 -683 -872
rect -625 -838 -465 -800
rect -625 -872 -609 -838
rect -481 -872 -465 -838
rect -625 -888 -465 -872
rect -407 -838 -247 -800
rect -407 -872 -391 -838
rect -263 -872 -247 -838
rect -407 -888 -247 -872
rect -189 -838 -29 -800
rect -189 -872 -173 -838
rect -45 -872 -29 -838
rect -189 -888 -29 -872
rect 29 -838 189 -800
rect 29 -872 45 -838
rect 173 -872 189 -838
rect 29 -888 189 -872
rect 247 -838 407 -800
rect 247 -872 263 -838
rect 391 -872 407 -838
rect 247 -888 407 -872
rect 465 -838 625 -800
rect 465 -872 481 -838
rect 609 -872 625 -838
rect 465 -888 625 -872
rect 683 -838 843 -800
rect 683 -872 699 -838
rect 827 -872 843 -838
rect 683 -888 843 -872
rect 901 -838 1061 -800
rect 901 -872 917 -838
rect 1045 -872 1061 -838
rect 901 -888 1061 -872
rect 1119 -838 1279 -800
rect 1119 -872 1135 -838
rect 1263 -872 1279 -838
rect 1119 -888 1279 -872
<< polycont >>
rect -1263 838 -1135 872
rect -1045 838 -917 872
rect -827 838 -699 872
rect -609 838 -481 872
rect -391 838 -263 872
rect -173 838 -45 872
rect 45 838 173 872
rect 263 838 391 872
rect 481 838 609 872
rect 699 838 827 872
rect 917 838 1045 872
rect 1135 838 1263 872
rect -1263 -872 -1135 -838
rect -1045 -872 -917 -838
rect -827 -872 -699 -838
rect -609 -872 -481 -838
rect -391 -872 -263 -838
rect -173 -872 -45 -838
rect 45 -872 173 -838
rect 263 -872 391 -838
rect 481 -872 609 -838
rect 699 -872 827 -838
rect 917 -872 1045 -838
rect 1135 -872 1263 -838
<< locali >>
rect -1459 976 -1363 1010
rect 1363 976 1459 1010
rect -1459 914 -1425 976
rect 1425 914 1459 976
rect -1279 838 -1263 872
rect -1135 838 -1119 872
rect -1061 838 -1045 872
rect -917 838 -901 872
rect -843 838 -827 872
rect -699 838 -683 872
rect -625 838 -609 872
rect -481 838 -465 872
rect -407 838 -391 872
rect -263 838 -247 872
rect -189 838 -173 872
rect -45 838 -29 872
rect 29 838 45 872
rect 173 838 189 872
rect 247 838 263 872
rect 391 838 407 872
rect 465 838 481 872
rect 609 838 625 872
rect 683 838 699 872
rect 827 838 843 872
rect 901 838 917 872
rect 1045 838 1061 872
rect 1119 838 1135 872
rect 1263 838 1279 872
rect -1325 788 -1291 804
rect -1325 -804 -1291 -788
rect -1107 788 -1073 804
rect -1107 -804 -1073 -788
rect -889 788 -855 804
rect -889 -804 -855 -788
rect -671 788 -637 804
rect -671 -804 -637 -788
rect -453 788 -419 804
rect -453 -804 -419 -788
rect -235 788 -201 804
rect -235 -804 -201 -788
rect -17 788 17 804
rect -17 -804 17 -788
rect 201 788 235 804
rect 201 -804 235 -788
rect 419 788 453 804
rect 419 -804 453 -788
rect 637 788 671 804
rect 637 -804 671 -788
rect 855 788 889 804
rect 855 -804 889 -788
rect 1073 788 1107 804
rect 1073 -804 1107 -788
rect 1291 788 1325 804
rect 1291 -804 1325 -788
rect -1279 -872 -1263 -838
rect -1135 -872 -1119 -838
rect -1061 -872 -1045 -838
rect -917 -872 -901 -838
rect -843 -872 -827 -838
rect -699 -872 -683 -838
rect -625 -872 -609 -838
rect -481 -872 -465 -838
rect -407 -872 -391 -838
rect -263 -872 -247 -838
rect -189 -872 -173 -838
rect -45 -872 -29 -838
rect 29 -872 45 -838
rect 173 -872 189 -838
rect 247 -872 263 -838
rect 391 -872 407 -838
rect 465 -872 481 -838
rect 609 -872 625 -838
rect 683 -872 699 -838
rect 827 -872 843 -838
rect 901 -872 917 -838
rect 1045 -872 1061 -838
rect 1119 -872 1135 -838
rect 1263 -872 1279 -838
rect -1459 -976 -1425 -914
rect 1425 -976 1459 -914
rect -1459 -1010 -1363 -976
rect 1363 -1010 1459 -976
<< viali >>
rect -1263 838 -1135 872
rect -1045 838 -917 872
rect -827 838 -699 872
rect -609 838 -481 872
rect -391 838 -263 872
rect -173 838 -45 872
rect 45 838 173 872
rect 263 838 391 872
rect 481 838 609 872
rect 699 838 827 872
rect 917 838 1045 872
rect 1135 838 1263 872
rect -1325 -788 -1291 788
rect -1107 -788 -1073 788
rect -889 -788 -855 788
rect -671 -788 -637 788
rect -453 -788 -419 788
rect -235 -788 -201 788
rect -17 -788 17 788
rect 201 -788 235 788
rect 419 -788 453 788
rect 637 -788 671 788
rect 855 -788 889 788
rect 1073 -788 1107 788
rect 1291 -788 1325 788
rect -1263 -872 -1135 -838
rect -1045 -872 -917 -838
rect -827 -872 -699 -838
rect -609 -872 -481 -838
rect -391 -872 -263 -838
rect -173 -872 -45 -838
rect 45 -872 173 -838
rect 263 -872 391 -838
rect 481 -872 609 -838
rect 699 -872 827 -838
rect 917 -872 1045 -838
rect 1135 -872 1263 -838
<< metal1 >>
rect -1275 872 -1123 878
rect -1275 838 -1263 872
rect -1135 838 -1123 872
rect -1275 832 -1123 838
rect -1057 872 -905 878
rect -1057 838 -1045 872
rect -917 838 -905 872
rect -1057 832 -905 838
rect -839 872 -687 878
rect -839 838 -827 872
rect -699 838 -687 872
rect -839 832 -687 838
rect -621 872 -469 878
rect -621 838 -609 872
rect -481 838 -469 872
rect -621 832 -469 838
rect -403 872 -251 878
rect -403 838 -391 872
rect -263 838 -251 872
rect -403 832 -251 838
rect -185 872 -33 878
rect -185 838 -173 872
rect -45 838 -33 872
rect -185 832 -33 838
rect 33 872 185 878
rect 33 838 45 872
rect 173 838 185 872
rect 33 832 185 838
rect 251 872 403 878
rect 251 838 263 872
rect 391 838 403 872
rect 251 832 403 838
rect 469 872 621 878
rect 469 838 481 872
rect 609 838 621 872
rect 469 832 621 838
rect 687 872 839 878
rect 687 838 699 872
rect 827 838 839 872
rect 687 832 839 838
rect 905 872 1057 878
rect 905 838 917 872
rect 1045 838 1057 872
rect 905 832 1057 838
rect 1123 872 1275 878
rect 1123 838 1135 872
rect 1263 838 1275 872
rect 1123 832 1275 838
rect -1331 788 -1285 800
rect -1331 -788 -1325 788
rect -1291 -788 -1285 788
rect -1331 -800 -1285 -788
rect -1113 788 -1067 800
rect -1113 -788 -1107 788
rect -1073 -788 -1067 788
rect -1113 -800 -1067 -788
rect -895 788 -849 800
rect -895 -788 -889 788
rect -855 -788 -849 788
rect -895 -800 -849 -788
rect -677 788 -631 800
rect -677 -788 -671 788
rect -637 -788 -631 788
rect -677 -800 -631 -788
rect -459 788 -413 800
rect -459 -788 -453 788
rect -419 -788 -413 788
rect -459 -800 -413 -788
rect -241 788 -195 800
rect -241 -788 -235 788
rect -201 -788 -195 788
rect -241 -800 -195 -788
rect -23 788 23 800
rect -23 -788 -17 788
rect 17 -788 23 788
rect -23 -800 23 -788
rect 195 788 241 800
rect 195 -788 201 788
rect 235 -788 241 788
rect 195 -800 241 -788
rect 413 788 459 800
rect 413 -788 419 788
rect 453 -788 459 788
rect 413 -800 459 -788
rect 631 788 677 800
rect 631 -788 637 788
rect 671 -788 677 788
rect 631 -800 677 -788
rect 849 788 895 800
rect 849 -788 855 788
rect 889 -788 895 788
rect 849 -800 895 -788
rect 1067 788 1113 800
rect 1067 -788 1073 788
rect 1107 -788 1113 788
rect 1067 -800 1113 -788
rect 1285 788 1331 800
rect 1285 -788 1291 788
rect 1325 -788 1331 788
rect 1285 -800 1331 -788
rect -1275 -838 -1123 -832
rect -1275 -872 -1263 -838
rect -1135 -872 -1123 -838
rect -1275 -878 -1123 -872
rect -1057 -838 -905 -832
rect -1057 -872 -1045 -838
rect -917 -872 -905 -838
rect -1057 -878 -905 -872
rect -839 -838 -687 -832
rect -839 -872 -827 -838
rect -699 -872 -687 -838
rect -839 -878 -687 -872
rect -621 -838 -469 -832
rect -621 -872 -609 -838
rect -481 -872 -469 -838
rect -621 -878 -469 -872
rect -403 -838 -251 -832
rect -403 -872 -391 -838
rect -263 -872 -251 -838
rect -403 -878 -251 -872
rect -185 -838 -33 -832
rect -185 -872 -173 -838
rect -45 -872 -33 -838
rect -185 -878 -33 -872
rect 33 -838 185 -832
rect 33 -872 45 -838
rect 173 -872 185 -838
rect 33 -878 185 -872
rect 251 -838 403 -832
rect 251 -872 263 -838
rect 391 -872 403 -838
rect 251 -878 403 -872
rect 469 -838 621 -832
rect 469 -872 481 -838
rect 609 -872 621 -838
rect 469 -878 621 -872
rect 687 -838 839 -832
rect 687 -872 699 -838
rect 827 -872 839 -838
rect 687 -878 839 -872
rect 905 -838 1057 -832
rect 905 -872 917 -838
rect 1045 -872 1057 -838
rect 905 -878 1057 -872
rect 1123 -838 1275 -832
rect 1123 -872 1135 -838
rect 1263 -872 1275 -838
rect 1123 -878 1275 -872
<< properties >>
string FIXED_BBOX -1442 -993 1442 993
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 8 l 0.8 m 1 nf 12 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
