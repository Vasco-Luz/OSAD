magic
tech sky130A
magscale 1 2
timestamp 1740407780
<< error_p >>
rect -353 548 353 552
rect -353 -480 -323 548
rect -287 482 287 486
rect -287 -414 -257 482
rect 257 -414 287 482
rect 323 -480 353 548
<< nwell >>
rect -323 -514 323 548
<< mvpmos >>
rect -229 -414 -29 486
rect 29 -414 229 486
<< mvpdiff >>
rect -287 474 -229 486
rect -287 -402 -275 474
rect -241 -402 -229 474
rect -287 -414 -229 -402
rect -29 474 29 486
rect -29 -402 -17 474
rect 17 -402 29 474
rect -29 -414 29 -402
rect 229 474 287 486
rect 229 -402 241 474
rect 275 -402 287 474
rect 229 -414 287 -402
<< mvpdiffc >>
rect -275 -402 -241 474
rect -17 -402 17 474
rect 241 -402 275 474
<< poly >>
rect -229 486 -29 512
rect 29 486 229 512
rect -229 -461 -29 -414
rect -229 -495 -213 -461
rect -45 -495 -29 -461
rect -229 -511 -29 -495
rect 29 -461 229 -414
rect 29 -495 45 -461
rect 213 -495 229 -461
rect 29 -511 229 -495
<< polycont >>
rect -213 -495 -45 -461
rect 45 -495 213 -461
<< locali >>
rect -275 474 -241 490
rect -275 -418 -241 -402
rect -17 474 17 490
rect -17 -418 17 -402
rect 241 474 275 490
rect 241 -418 275 -402
rect -229 -495 -213 -461
rect -45 -495 -29 -461
rect 29 -495 45 -461
rect 213 -495 229 -461
<< viali >>
rect -275 -402 -241 474
rect -17 -402 17 474
rect 241 -402 275 474
rect -196 -495 -62 -461
rect 62 -495 196 -461
<< metal1 >>
rect -275 486 -241 596
rect -17 486 17 622
rect 241 486 275 618
rect -281 474 -235 486
rect -281 -402 -275 474
rect -241 -402 -235 474
rect -281 -414 -235 -402
rect -23 474 23 486
rect -23 -402 -17 474
rect 17 -402 23 474
rect -23 -414 23 -402
rect 235 474 281 486
rect 235 -402 241 474
rect 275 -402 281 474
rect 235 -414 281 -402
rect -208 -461 -50 -455
rect -208 -495 -196 -461
rect -62 -495 -50 -461
rect -208 -501 -50 -495
rect 50 -461 208 -455
rect 50 -495 62 -461
rect 196 -495 208 -461
rect 50 -501 208 -495
rect -93 -738 -61 -501
rect 165 -736 197 -501
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 4.5 l 1 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 80 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 80 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
