magic
tech sky130A
magscale 1 2
timestamp 1730736629
<< nmos >>
rect -600 708 0 1108
rect 58 708 658 1108
rect 716 708 1316 1108
rect 1374 708 1974 1108
rect 2032 708 2632 1108
rect 2690 708 3290 1108
rect 3348 708 3948 1108
rect 4006 708 4606 1108
rect 4664 708 5264 1108
rect 5322 708 5922 1108
rect 5980 708 6580 1108
rect 6638 708 7238 1108
rect 7296 708 7896 1108
rect 7954 708 8554 1108
<< ndiff >>
rect -658 1096 -600 1108
rect -658 720 -646 1096
rect -612 720 -600 1096
rect -658 708 -600 720
rect 0 1096 58 1108
rect 0 720 12 1096
rect 46 720 58 1096
rect 0 708 58 720
rect 658 1096 716 1108
rect 658 720 670 1096
rect 704 720 716 1096
rect 658 708 716 720
rect 1316 1096 1374 1108
rect 1316 720 1328 1096
rect 1362 720 1374 1096
rect 1316 708 1374 720
rect 1974 1096 2032 1108
rect 1974 720 1986 1096
rect 2020 720 2032 1096
rect 1974 708 2032 720
rect 2632 1096 2690 1108
rect 2632 720 2644 1096
rect 2678 720 2690 1096
rect 2632 708 2690 720
rect 3290 1096 3348 1108
rect 3290 720 3302 1096
rect 3336 720 3348 1096
rect 3290 708 3348 720
rect 3948 1096 4006 1108
rect 3948 720 3960 1096
rect 3994 720 4006 1096
rect 3948 708 4006 720
rect 4606 1096 4664 1108
rect 4606 720 4618 1096
rect 4652 720 4664 1096
rect 4606 708 4664 720
rect 5264 1096 5322 1108
rect 5264 720 5276 1096
rect 5310 720 5322 1096
rect 5264 708 5322 720
rect 5922 1096 5980 1108
rect 5922 720 5934 1096
rect 5968 720 5980 1096
rect 5922 708 5980 720
rect 6580 1096 6638 1108
rect 6580 720 6592 1096
rect 6626 720 6638 1096
rect 6580 708 6638 720
rect 7238 1096 7296 1108
rect 7238 720 7250 1096
rect 7284 720 7296 1096
rect 7238 708 7296 720
rect 7896 1096 7954 1108
rect 7896 720 7908 1096
rect 7942 720 7954 1096
rect 7896 708 7954 720
rect 8554 1096 8612 1108
rect 8554 720 8566 1096
rect 8600 720 8612 1096
rect 8554 708 8612 720
<< ndiffc >>
rect -646 720 -612 1096
rect 12 720 46 1096
rect 670 720 704 1096
rect 1328 720 1362 1096
rect 1986 720 2020 1096
rect 2644 720 2678 1096
rect 3302 720 3336 1096
rect 3960 720 3994 1096
rect 4618 720 4652 1096
rect 5276 720 5310 1096
rect 5934 720 5968 1096
rect 6592 720 6626 1096
rect 7250 720 7284 1096
rect 7908 720 7942 1096
rect 8566 720 8600 1096
<< psubdiff >>
rect -809 1303 -749 1337
rect 8723 1303 8783 1337
rect -809 1277 -775 1303
rect 8749 1277 8783 1303
rect -809 -137 -775 -111
rect 8749 -137 8783 -111
rect -809 -171 -749 -137
rect 8723 -171 8783 -137
<< psubdiffcont >>
rect -749 1303 8723 1337
rect -809 -111 -775 1277
rect 8749 -111 8783 1277
rect -749 -171 8723 -137
<< poly >>
rect -600 1108 0 1134
rect 58 1108 658 1134
rect 716 1108 1316 1134
rect 1374 1108 1974 1134
rect 2032 1108 2632 1134
rect 2690 1108 3290 1134
rect 3348 1108 3948 1134
rect 4006 1108 4606 1134
rect 4664 1108 5264 1134
rect 5322 1108 5922 1134
rect 5980 1108 6580 1134
rect 6638 1108 7238 1134
rect 7296 1108 7896 1134
rect 7954 1108 8554 1134
rect -600 682 0 708
rect 58 682 658 708
rect 716 682 1316 708
rect 1374 682 1974 708
rect 2032 682 2632 708
rect 2690 682 3290 708
rect 3348 682 3948 708
rect 4006 682 4606 708
rect 4664 682 5264 708
rect 5322 682 5922 708
rect 5980 682 6580 708
rect 6638 682 7238 708
rect 7296 682 7896 708
rect 7954 682 8554 708
<< locali >>
rect -809 1303 -749 1337
rect 8723 1303 8783 1337
rect -809 1277 -775 1303
rect 8749 1277 8783 1303
rect -646 1096 -612 1112
rect -646 704 -612 720
rect 12 1096 46 1112
rect 12 704 46 720
rect 670 1096 704 1112
rect 670 704 704 720
rect 1328 1096 1362 1112
rect 1328 704 1362 720
rect 1986 1096 2020 1112
rect 1986 704 2020 720
rect 2644 1096 2678 1112
rect 2644 704 2678 720
rect 3302 1096 3336 1112
rect 3302 704 3336 720
rect 3960 1096 3994 1112
rect 3960 704 3994 720
rect 4618 1096 4652 1112
rect 4618 704 4652 720
rect 5276 1096 5310 1112
rect 5276 704 5310 720
rect 5934 1096 5968 1112
rect 5934 704 5968 720
rect 6592 1096 6626 1112
rect 6592 704 6626 720
rect 7250 1096 7284 1112
rect 7250 704 7284 720
rect 7908 1096 7942 1112
rect 7908 704 7942 720
rect 8566 1096 8600 1112
rect 8566 704 8600 720
rect -809 -137 -775 -111
rect 8749 -137 8783 -111
rect -809 -171 -749 -137
rect 8723 -171 8783 -137
<< viali >>
rect -646 720 -612 1096
rect 12 720 46 1096
rect 670 720 704 1096
rect 1328 720 1362 1096
rect 1986 720 2020 1096
rect 2644 720 2678 1096
rect 3302 720 3336 1096
rect 3960 720 3994 1096
rect 4618 720 4652 1096
rect 5276 720 5310 1096
rect 5934 720 5968 1096
rect 6592 720 6626 1096
rect 7250 720 7284 1096
rect 7908 720 7942 1096
rect 8566 720 8600 1096
<< metal1 >>
rect -652 1096 -606 1108
rect -652 720 -646 1096
rect -612 720 -606 1096
rect -652 708 -606 720
rect 6 1096 52 1108
rect 6 720 12 1096
rect 46 720 52 1096
rect 6 708 52 720
rect 664 1096 710 1108
rect 664 720 670 1096
rect 704 720 710 1096
rect 664 708 710 720
rect 1322 1096 1368 1108
rect 1322 720 1328 1096
rect 1362 720 1368 1096
rect 1322 708 1368 720
rect 1980 1096 2026 1108
rect 1980 720 1986 1096
rect 2020 720 2026 1096
rect 1980 708 2026 720
rect 2638 1096 2684 1108
rect 2638 720 2644 1096
rect 2678 720 2684 1096
rect 2638 708 2684 720
rect 3296 1096 3342 1108
rect 3296 720 3302 1096
rect 3336 720 3342 1096
rect 3296 708 3342 720
rect 3954 1096 4000 1108
rect 3954 720 3960 1096
rect 3994 720 4000 1096
rect 3954 708 4000 720
rect 4612 1096 4658 1108
rect 4612 720 4618 1096
rect 4652 720 4658 1096
rect 4612 708 4658 720
rect 5270 1096 5316 1108
rect 5270 720 5276 1096
rect 5310 720 5316 1096
rect 5270 708 5316 720
rect 5928 1096 5974 1108
rect 5928 720 5934 1096
rect 5968 720 5974 1096
rect 5928 708 5974 720
rect 6586 1096 6632 1108
rect 6586 720 6592 1096
rect 6626 720 6632 1096
rect 6586 708 6632 720
rect 7244 1096 7290 1108
rect 7244 720 7250 1096
rect 7284 720 7290 1096
rect 7244 708 7290 720
rect 7902 1096 7948 1108
rect 7902 720 7908 1096
rect 7942 720 7948 1096
rect 7902 708 7948 720
rect 8560 1096 8606 1108
rect 8560 720 8566 1096
rect 8600 720 8606 1096
rect 8560 708 8606 720
use sky130_fd_pr__nfet_01v8_3TJNGK  sky130_fd_pr__nfet_01v8_3TJNGK_0
timestamp 1730731387
transform 1 0 2990 0 1 226
box -358 -226 358 226
use sky130_fd_pr__nfet_01v8_3TJNGK  sky130_fd_pr__nfet_01v8_3TJNGK_1
timestamp 1730731387
transform 1 0 4306 0 1 226
box -358 -226 358 226
use sky130_fd_pr__nfet_01v8_3TJNGK  sky130_fd_pr__nfet_01v8_3TJNGK_2
timestamp 1730731387
transform 1 0 358 0 1 226
box -358 -226 358 226
use sky130_fd_pr__nfet_01v8_3TJNGK  sky130_fd_pr__nfet_01v8_3TJNGK_3
timestamp 1730731387
transform 1 0 1016 0 1 226
box -358 -226 358 226
use sky130_fd_pr__nfet_01v8_3TJNGK  sky130_fd_pr__nfet_01v8_3TJNGK_4
timestamp 1730731387
transform 1 0 -300 0 1 226
box -358 -226 358 226
use sky130_fd_pr__nfet_01v8_3TJNGK  sky130_fd_pr__nfet_01v8_3TJNGK_5
timestamp 1730731387
transform 1 0 1674 0 1 226
box -358 -226 358 226
use sky130_fd_pr__nfet_01v8_3TJNGK  sky130_fd_pr__nfet_01v8_3TJNGK_6
timestamp 1730731387
transform 1 0 2332 0 1 226
box -358 -226 358 226
use sky130_fd_pr__nfet_01v8_3TJNGK  sky130_fd_pr__nfet_01v8_3TJNGK_7
timestamp 1730731387
transform 1 0 5622 0 1 226
box -358 -226 358 226
use sky130_fd_pr__nfet_01v8_3TJNGK  sky130_fd_pr__nfet_01v8_3TJNGK_8
timestamp 1730731387
transform 1 0 3648 0 1 226
box -358 -226 358 226
use sky130_fd_pr__nfet_01v8_3TJNGK  sky130_fd_pr__nfet_01v8_3TJNGK_9
timestamp 1730731387
transform 1 0 4964 0 1 226
box -358 -226 358 226
use sky130_fd_pr__nfet_01v8_3TJNGK *sky130_fd_pr__nfet_01v8_3TJNGK_10
timestamp 1730731387
transform 1 0 8254 0 1 226
box -358 -226 358 226
use sky130_fd_pr__nfet_01v8_3TJNGK  sky130_fd_pr__nfet_01v8_3TJNGK_11
timestamp 1730731387
transform 1 0 6280 0 1 226
box -358 -226 358 226
use sky130_fd_pr__nfet_01v8_3TJNGK  sky130_fd_pr__nfet_01v8_3TJNGK_12
timestamp 1730731387
transform 1 0 6938 0 1 226
box -358 -226 358 226
use sky130_fd_pr__nfet_01v8_3TJNGK *sky130_fd_pr__nfet_01v8_3TJNGK_14
timestamp 1730731387
transform 1 0 7596 0 1 226
box -358 -226 358 226
<< labels >>
flabel nmos 6748 778 7128 1040 0 FreeSans 800 0 0 0 M3
flabel nmos 6098 774 6460 1044 0 FreeSans 800 0 0 0 Dummy
flabel nmos 7412 750 7746 1044 0 FreeSans 800 0 0 0 M3
flabel nmos 8126 780 8460 1074 0 FreeSans 800 0 0 0 Dummy
flabel nmos -458 744 -128 994 0 FreeSans 800 0 0 0 dummy
flabel nmos 224 826 590 1006 0 FreeSans 800 0 0 0 M3
flabel nmos 830 814 1176 1014 0 FreeSans 800 0 0 0 M3
flabel nmos 1452 782 1844 1036 0 FreeSans 800 0 0 0 Dummy
flabel nmos 2142 766 2534 1020 0 FreeSans 800 0 0 0 Dummy
flabel nmos 2762 780 3130 1028 0 FreeSans 800 0 0 0 M4
flabel nmos 3500 808 3742 970 0 FreeSans 800 0 0 0 M4
flabel nmos 4108 812 4400 970 0 FreeSans 800 0 0 0 M4
flabel nmos 4808 808 5060 968 0 FreeSans 800 0 0 0 M4
flabel nmos 5418 762 5786 1054 0 FreeSans 800 0 0 0 Dummy
flabel space 8126 98 8460 392 0 FreeSans 800 0 0 0 Dummy
flabel space 7412 68 7746 362 0 FreeSans 800 0 0 0 M3
flabel space 6748 96 7128 358 0 FreeSans 800 0 0 0 M3
flabel space 6098 92 6460 362 0 FreeSans 800 0 0 0 Dummy
flabel space 5418 80 5786 372 0 FreeSans 800 0 0 0 Dummy
flabel space 4808 126 5060 286 0 FreeSans 800 0 0 0 M4
flabel space 4108 130 4400 288 0 FreeSans 800 0 0 0 M4
flabel space 3500 126 3742 288 0 FreeSans 800 0 0 0 M4
flabel space 2762 98 3130 346 0 FreeSans 800 0 0 0 M4
flabel space 2142 84 2534 338 0 FreeSans 800 0 0 0 Dummy
flabel space 1452 100 1844 354 0 FreeSans 800 0 0 0 Dummy
flabel space 830 132 1176 332 0 FreeSans 800 0 0 0 M3
flabel space 224 144 590 324 0 FreeSans 800 0 0 0 M3
flabel space -458 62 -128 312 0 FreeSans 800 0 0 0 dummy
<< end >>
