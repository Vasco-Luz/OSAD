** sch_path: /home/vasco/Desktop/OSAD/my_ip/testbenches_sky/transcondutance_cell/test.sch
**.subckt test
V1 VDD GND VDD
V2 VSS GND VSS
XM2 net4 net3 net2 net2 sky130_fd_pr__pfet_g5v0d10v5 L=2.8 W=2.7 nf=4 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=3 m=3
XM1 net3 net3 net1 net1 sky130_fd_pr__pfet_g5v0d10v5 L=2.8 W=2.7 nf=4 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=3 m=3
XM4 net4 net4 net5 VSS sky130_fd_pr__nfet_g5v0d10v5 L=2.8 W=2.7 nf=8 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
XM3 net3 net4 net6 VSS sky130_fd_pr__nfet_g5v0d10v5 L=2.8 W=2.7 nf=8 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
XM5 net6 net5 net7 VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=1.5 nf=6 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=16 m=16
XR6 VSS net7 VSS sky130_fd_pr__res_high_po_0p35 L=2.5 mult=1 m=1
Vmeas VDD net1 0
.save i(vmeas)
Vmeas1 VDD net2 0
.save i(vmeas1)
XM6 net5 net5 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=1.5 nf=6 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4
**** begin user architecture code
.lib /home/vasco/PDK/sky130A/libs.tech/combined/sky130.lib.spice tt
.Temp 27
.param VDD = 5
.param VSS = 0
.control
save all
dc Temp -40 125 1
plot i(Vmeas) i(Vmeas1)
wrdata transimpedance.csv i(Vmeas) i(Vmeas1)
.endc
**** end user architecture code
**.ends
.GLOBAL GND
.end