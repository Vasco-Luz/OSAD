magic
tech sky130A
magscale 1 2
timestamp 1730740146
<< poly >>
rect 213 1404 813 1424
rect 213 1370 412 1404
rect 632 1370 813 1404
rect 213 1305 813 1370
rect 871 1404 1471 1424
rect 871 1370 1070 1404
rect 1290 1370 1471 1404
rect 871 1305 1471 1370
rect 1529 1404 2129 1424
rect 1529 1370 1728 1404
rect 1948 1370 2129 1404
rect 1529 1305 2129 1370
rect 2187 1404 2787 1424
rect 2187 1370 2386 1404
rect 2606 1370 2787 1404
rect 2187 1305 2787 1370
rect 2845 1404 3445 1424
rect 2845 1370 3044 1404
rect 3264 1370 3445 1404
rect 2845 1305 3445 1370
rect 3503 1404 4103 1424
rect 3503 1370 3702 1404
rect 3922 1370 4103 1404
rect 3503 1305 4103 1370
rect 4161 1404 4761 1424
rect 4161 1370 4360 1404
rect 4580 1370 4761 1404
rect 4161 1305 4761 1370
rect 4819 1423 5419 1443
rect 4819 1389 5018 1423
rect 5238 1389 5419 1423
rect 4819 1305 5419 1389
rect 5477 1423 6077 1443
rect 5477 1389 5676 1423
rect 5896 1389 6077 1423
rect 5477 1305 6077 1389
rect 6135 1423 6735 1443
rect 6135 1389 6334 1423
rect 6554 1389 6735 1423
rect 6135 1305 6735 1389
rect 6793 1423 7393 1443
rect 6793 1389 6992 1423
rect 7212 1389 7393 1423
rect 6793 1305 7393 1389
rect 7451 1423 8051 1443
rect 7451 1389 7650 1423
rect 7870 1389 8051 1423
rect 7451 1305 8051 1389
rect 8109 1423 8709 1443
rect 8109 1389 8308 1423
rect 8528 1389 8709 1423
rect 8109 1305 8709 1389
rect 8767 1423 9367 1443
rect 8767 1389 8966 1423
rect 9186 1389 9367 1423
rect 8767 1305 9367 1389
rect 4819 716 5419 736
rect 4819 682 5018 716
rect 5238 682 5419 716
rect 4819 623 5419 682
rect 5477 716 6077 736
rect 5477 682 5676 716
rect 5896 682 6077 716
rect 5477 623 6077 682
rect 6135 716 6735 736
rect 6135 682 6334 716
rect 6554 682 6735 716
rect 6135 623 6735 682
rect 6793 716 7393 736
rect 6793 682 6992 716
rect 7212 682 7393 716
rect 6793 623 7393 682
rect 7451 716 8051 736
rect 7451 682 7650 716
rect 7870 682 8051 716
rect 7451 623 8051 682
rect 8109 716 8709 736
rect 8109 682 8308 716
rect 8528 682 8709 716
rect 8109 623 8709 682
rect 8767 716 9367 736
rect 8767 682 8966 716
rect 9186 682 9367 716
rect 8767 623 9367 682
<< polycont >>
rect 412 1370 632 1404
rect 1070 1370 1290 1404
rect 1728 1370 1948 1404
rect 2386 1370 2606 1404
rect 3044 1370 3264 1404
rect 3702 1370 3922 1404
rect 4360 1370 4580 1404
rect 5018 1389 5238 1423
rect 5676 1389 5896 1423
rect 6334 1389 6554 1423
rect 6992 1389 7212 1423
rect 7650 1389 7870 1423
rect 8308 1389 8528 1423
rect 8966 1389 9186 1423
rect 5018 682 5238 716
rect 5676 682 5896 716
rect 6334 682 6554 716
rect 6992 682 7212 716
rect 7650 682 7870 716
rect 8308 682 8528 716
rect 8966 682 9186 716
<< locali >>
rect 166 4 202 1484
rect 5002 1423 5254 1439
rect 396 1404 648 1420
rect 396 1370 412 1404
rect 632 1370 648 1404
rect 396 1354 648 1370
rect 1054 1404 1306 1420
rect 1054 1370 1070 1404
rect 1290 1370 1306 1404
rect 1054 1354 1306 1370
rect 1712 1404 1964 1420
rect 1712 1370 1728 1404
rect 1948 1370 1964 1404
rect 1712 1354 1964 1370
rect 2370 1404 2622 1420
rect 2370 1370 2386 1404
rect 2606 1370 2622 1404
rect 2370 1354 2622 1370
rect 3028 1404 3280 1420
rect 3028 1370 3044 1404
rect 3264 1370 3280 1404
rect 3028 1354 3280 1370
rect 3686 1404 3938 1420
rect 3686 1370 3702 1404
rect 3922 1370 3938 1404
rect 3686 1354 3938 1370
rect 4344 1404 4596 1420
rect 4344 1370 4360 1404
rect 4580 1370 4596 1404
rect 5002 1389 5018 1423
rect 5238 1389 5254 1423
rect 5002 1373 5254 1389
rect 5660 1423 5912 1439
rect 5660 1389 5676 1423
rect 5896 1389 5912 1423
rect 5660 1373 5912 1389
rect 6318 1423 6570 1439
rect 6318 1389 6334 1423
rect 6554 1389 6570 1423
rect 6318 1373 6570 1389
rect 6976 1423 7228 1439
rect 6976 1389 6992 1423
rect 7212 1389 7228 1423
rect 6976 1373 7228 1389
rect 7634 1423 7886 1439
rect 7634 1389 7650 1423
rect 7870 1389 7886 1423
rect 7634 1373 7886 1389
rect 8292 1423 8544 1439
rect 8292 1389 8308 1423
rect 8528 1389 8544 1423
rect 8292 1373 8544 1389
rect 8950 1423 9202 1439
rect 8950 1389 8966 1423
rect 9186 1389 9202 1423
rect 8950 1373 9202 1389
rect 4344 1354 4596 1370
rect 5002 716 5254 732
rect 5002 682 5018 716
rect 5238 682 5254 716
rect 5002 666 5254 682
rect 5660 716 5912 732
rect 5660 682 5676 716
rect 5896 682 5912 716
rect 5660 666 5912 682
rect 6318 716 6570 732
rect 6318 682 6334 716
rect 6554 682 6570 716
rect 6318 666 6570 682
rect 6976 716 7228 732
rect 6976 682 6992 716
rect 7212 682 7228 716
rect 6976 666 7228 682
rect 7634 716 7886 732
rect 7634 682 7650 716
rect 7870 682 7886 716
rect 7634 666 7886 682
rect 8292 716 8544 732
rect 8292 682 8308 716
rect 8528 682 8544 716
rect 8292 666 8544 682
rect 8950 716 9202 732
rect 8950 682 8966 716
rect 9186 682 9202 716
rect 8950 666 9202 682
<< viali >>
rect 412 1370 632 1404
rect 1070 1370 1290 1404
rect 1728 1370 1948 1404
rect 2386 1370 2606 1404
rect 3044 1370 3264 1404
rect 3702 1370 3922 1404
rect 4360 1370 4580 1404
rect 5018 1389 5238 1423
rect 5676 1389 5896 1423
rect 6334 1389 6554 1423
rect 6992 1389 7212 1423
rect 7650 1389 7870 1423
rect 8308 1389 8528 1423
rect 8966 1389 9186 1423
rect 5018 682 5238 716
rect 5676 682 5896 716
rect 6334 682 6554 716
rect 6992 682 7212 716
rect 7650 682 7870 716
rect 8308 682 8528 716
rect 8966 682 9186 716
<< metal1 >>
rect 5006 1423 5250 1435
rect 400 1404 644 1416
rect 400 1370 412 1404
rect 632 1370 644 1404
rect 400 1356 644 1370
rect 1058 1404 1302 1416
rect 1058 1370 1070 1404
rect 1290 1370 1302 1404
rect 1058 1356 1302 1370
rect 1716 1404 1960 1416
rect 1716 1370 1728 1404
rect 1948 1370 1960 1404
rect 1716 1356 1960 1370
rect 2374 1404 2618 1416
rect 2374 1370 2386 1404
rect 2606 1370 2618 1404
rect 2374 1356 2618 1370
rect 3032 1404 3276 1416
rect 3032 1370 3044 1404
rect 3264 1370 3276 1404
rect 3032 1356 3276 1370
rect 3690 1404 3934 1416
rect 3690 1370 3702 1404
rect 3922 1370 3934 1404
rect 3690 1356 3934 1370
rect 4348 1404 4592 1416
rect 4348 1370 4360 1404
rect 4580 1370 4592 1404
rect 5006 1389 5018 1423
rect 5238 1389 5250 1423
rect 5006 1375 5250 1389
rect 5664 1423 5908 1435
rect 5664 1389 5676 1423
rect 5896 1389 5908 1423
rect 5664 1375 5908 1389
rect 6322 1423 6566 1435
rect 6322 1389 6334 1423
rect 6554 1389 6566 1423
rect 6322 1375 6566 1389
rect 6980 1423 7224 1435
rect 6980 1389 6992 1423
rect 7212 1389 7224 1423
rect 6980 1375 7224 1389
rect 7638 1423 7882 1435
rect 7638 1389 7650 1423
rect 7870 1389 7882 1423
rect 7638 1375 7882 1389
rect 8296 1423 8540 1435
rect 8296 1389 8308 1423
rect 8528 1389 8540 1423
rect 8296 1375 8540 1389
rect 8954 1423 9198 1435
rect 8954 1389 8966 1423
rect 9186 1389 9198 1423
rect 8954 1375 9198 1389
rect 4348 1356 4592 1370
rect 5006 716 5250 728
rect 5006 682 5018 716
rect 5238 682 5250 716
rect 5006 668 5250 682
rect 5664 716 5908 728
rect 5664 682 5676 716
rect 5896 682 5908 716
rect 5664 668 5908 682
rect 6322 716 6566 728
rect 6322 682 6334 716
rect 6554 682 6566 716
rect 6322 668 6566 682
rect 6980 716 7224 728
rect 6980 682 6992 716
rect 7212 682 7224 716
rect 6980 668 7224 682
rect 7638 716 7882 728
rect 7638 682 7650 716
rect 7870 682 7882 716
rect 7638 668 7882 682
rect 8296 716 8540 728
rect 8296 682 8308 716
rect 8528 682 8540 716
rect 8296 668 8540 682
rect 8954 716 9198 728
rect 8954 682 8966 716
rect 9186 682 9198 716
rect 8954 668 9198 682
use NMOS_higher_first  NMOS_higher_first_0
timestamp 1730736629
transform 1 0 813 0 1 171
box -809 -171 8783 1337
use NMOS_UPPER_contact_gate  NMOS_UPPER_contact_gate_0
timestamp 1730737099
transform 1 0 3950 0 1 27
box 211 596 811 690
use NMOS_UPPER_contact_gate  NMOS_UPPER_contact_gate_1
timestamp 1730737099
transform 1 0 2 0 1 27
box 211 596 811 690
use NMOS_UPPER_contact_gate  NMOS_UPPER_contact_gate_2
timestamp 1730737099
transform 1 0 660 0 1 27
box 211 596 811 690
use NMOS_UPPER_contact_gate  NMOS_UPPER_contact_gate_3
timestamp 1730737099
transform 1 0 1318 0 1 27
box 211 596 811 690
use NMOS_UPPER_contact_gate  NMOS_UPPER_contact_gate_4
timestamp 1730737099
transform 1 0 1976 0 1 27
box 211 596 811 690
use NMOS_UPPER_contact_gate  NMOS_UPPER_contact_gate_5
timestamp 1730737099
transform 1 0 2634 0 1 27
box 211 596 811 690
use NMOS_UPPER_contact_gate  NMOS_UPPER_contact_gate_6
timestamp 1730737099
transform 1 0 3292 0 1 27
box 211 596 811 690
<< end >>
