magic
tech sky130A
magscale 1 2
timestamp 1740407780
<< error_p >>
rect -611 548 611 552
rect -611 -480 -581 548
rect -545 482 545 486
rect -545 -414 -515 482
rect 515 -414 545 482
rect 581 -480 611 548
<< nwell >>
rect -581 -514 581 548
<< mvpmos >>
rect -487 -414 -287 486
rect -229 -414 -29 486
rect 29 -414 229 486
rect 287 -414 487 486
<< mvpdiff >>
rect -545 474 -487 486
rect -545 -402 -533 474
rect -499 -402 -487 474
rect -545 -414 -487 -402
rect -287 474 -229 486
rect -287 -402 -275 474
rect -241 -402 -229 474
rect -287 -414 -229 -402
rect -29 474 29 486
rect -29 -402 -17 474
rect 17 -402 29 474
rect -29 -414 29 -402
rect 229 474 287 486
rect 229 -402 241 474
rect 275 -402 287 474
rect 229 -414 287 -402
rect 487 474 545 486
rect 487 -402 499 474
rect 533 -402 545 474
rect 487 -414 545 -402
<< mvpdiffc >>
rect -533 -402 -499 474
rect -275 -402 -241 474
rect -17 -402 17 474
rect 241 -402 275 474
rect 499 -402 533 474
<< poly >>
rect -487 486 -287 512
rect -229 486 -29 512
rect 29 486 229 512
rect 287 486 487 512
rect -487 -461 -287 -414
rect -487 -495 -471 -461
rect -303 -495 -287 -461
rect -487 -511 -287 -495
rect -229 -461 -29 -414
rect -229 -495 -213 -461
rect -45 -495 -29 -461
rect -229 -511 -29 -495
rect 29 -461 229 -414
rect 29 -495 45 -461
rect 213 -495 229 -461
rect 29 -511 229 -495
rect 287 -461 487 -414
rect 287 -495 303 -461
rect 471 -495 487 -461
rect 287 -511 487 -495
<< polycont >>
rect -471 -495 -303 -461
rect -213 -495 -45 -461
rect 45 -495 213 -461
rect 303 -495 471 -461
<< locali >>
rect -533 474 -499 490
rect -533 -418 -499 -402
rect -275 474 -241 490
rect -275 -418 -241 -402
rect -17 474 17 490
rect -17 -418 17 -402
rect 241 474 275 490
rect 241 -418 275 -402
rect 499 474 533 490
rect 499 -418 533 -402
rect -487 -495 -471 -461
rect -303 -495 -287 -461
rect -229 -495 -213 -461
rect -45 -495 -29 -461
rect 29 -495 45 -461
rect 213 -495 229 -461
rect 287 -495 303 -461
rect 471 -495 487 -461
<< viali >>
rect -533 -402 -499 474
rect -275 -402 -241 474
rect -17 -402 17 474
rect 241 -402 275 474
rect 499 -402 533 474
rect -454 -495 -320 -461
rect -196 -495 -62 -461
rect 62 -495 196 -461
rect 320 -495 454 -461
<< metal1 >>
rect -539 474 -493 486
rect -539 -402 -533 474
rect -499 -402 -493 474
rect -539 -414 -493 -402
rect -281 474 -235 486
rect -281 -402 -275 474
rect -241 -402 -235 474
rect -281 -414 -235 -402
rect -23 474 23 486
rect -23 -402 -17 474
rect 17 -402 23 474
rect -23 -414 23 -402
rect 235 474 281 486
rect 235 -402 241 474
rect 275 -402 281 474
rect 235 -414 281 -402
rect 493 474 539 486
rect 493 -402 499 474
rect 533 -402 539 474
rect 493 -414 539 -402
rect -466 -461 -308 -455
rect -466 -495 -454 -461
rect -320 -495 -308 -461
rect -466 -501 -308 -495
rect -208 -461 -50 -455
rect -208 -495 -196 -461
rect -62 -495 -50 -461
rect -208 -501 -50 -495
rect 50 -461 208 -455
rect 50 -495 62 -461
rect 196 -495 208 -461
rect 50 -501 208 -495
rect 308 -461 466 -455
rect 308 -495 320 -461
rect 454 -495 466 -461
rect 308 -501 466 -495
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 4.5 l 1 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 80 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 80 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
