magic
tech sky130A
magscale 1 2
timestamp 1693698878
<< nwell >>
rect -1537 -697 1537 697
<< mvpmos >>
rect -1279 -400 -1119 400
rect -1061 -400 -901 400
rect -843 -400 -683 400
rect -625 -400 -465 400
rect -407 -400 -247 400
rect -189 -400 -29 400
rect 29 -400 189 400
rect 247 -400 407 400
rect 465 -400 625 400
rect 683 -400 843 400
rect 901 -400 1061 400
rect 1119 -400 1279 400
<< mvpdiff >>
rect -1337 388 -1279 400
rect -1337 -388 -1325 388
rect -1291 -388 -1279 388
rect -1337 -400 -1279 -388
rect -1119 388 -1061 400
rect -1119 -388 -1107 388
rect -1073 -388 -1061 388
rect -1119 -400 -1061 -388
rect -901 388 -843 400
rect -901 -388 -889 388
rect -855 -388 -843 388
rect -901 -400 -843 -388
rect -683 388 -625 400
rect -683 -388 -671 388
rect -637 -388 -625 388
rect -683 -400 -625 -388
rect -465 388 -407 400
rect -465 -388 -453 388
rect -419 -388 -407 388
rect -465 -400 -407 -388
rect -247 388 -189 400
rect -247 -388 -235 388
rect -201 -388 -189 388
rect -247 -400 -189 -388
rect -29 388 29 400
rect -29 -388 -17 388
rect 17 -388 29 388
rect -29 -400 29 -388
rect 189 388 247 400
rect 189 -388 201 388
rect 235 -388 247 388
rect 189 -400 247 -388
rect 407 388 465 400
rect 407 -388 419 388
rect 453 -388 465 388
rect 407 -400 465 -388
rect 625 388 683 400
rect 625 -388 637 388
rect 671 -388 683 388
rect 625 -400 683 -388
rect 843 388 901 400
rect 843 -388 855 388
rect 889 -388 901 388
rect 843 -400 901 -388
rect 1061 388 1119 400
rect 1061 -388 1073 388
rect 1107 -388 1119 388
rect 1061 -400 1119 -388
rect 1279 388 1337 400
rect 1279 -388 1291 388
rect 1325 -388 1337 388
rect 1279 -400 1337 -388
<< mvpdiffc >>
rect -1325 -388 -1291 388
rect -1107 -388 -1073 388
rect -889 -388 -855 388
rect -671 -388 -637 388
rect -453 -388 -419 388
rect -235 -388 -201 388
rect -17 -388 17 388
rect 201 -388 235 388
rect 419 -388 453 388
rect 637 -388 671 388
rect 855 -388 889 388
rect 1073 -388 1107 388
rect 1291 -388 1325 388
<< mvnsubdiff >>
rect -1471 619 1471 631
rect -1471 585 -1363 619
rect 1363 585 1471 619
rect -1471 573 1471 585
rect -1471 523 -1413 573
rect -1471 -523 -1459 523
rect -1425 -523 -1413 523
rect 1413 523 1471 573
rect -1471 -573 -1413 -523
rect 1413 -523 1425 523
rect 1459 -523 1471 523
rect 1413 -573 1471 -523
rect -1471 -585 1471 -573
rect -1471 -619 -1363 -585
rect 1363 -619 1471 -585
rect -1471 -631 1471 -619
<< mvnsubdiffcont >>
rect -1363 585 1363 619
rect -1459 -523 -1425 523
rect 1425 -523 1459 523
rect -1363 -619 1363 -585
<< poly >>
rect -1279 481 -1119 497
rect -1279 447 -1263 481
rect -1135 447 -1119 481
rect -1279 400 -1119 447
rect -1061 481 -901 497
rect -1061 447 -1045 481
rect -917 447 -901 481
rect -1061 400 -901 447
rect -843 481 -683 497
rect -843 447 -827 481
rect -699 447 -683 481
rect -843 400 -683 447
rect -625 481 -465 497
rect -625 447 -609 481
rect -481 447 -465 481
rect -625 400 -465 447
rect -407 481 -247 497
rect -407 447 -391 481
rect -263 447 -247 481
rect -407 400 -247 447
rect -189 481 -29 497
rect -189 447 -173 481
rect -45 447 -29 481
rect -189 400 -29 447
rect 29 481 189 497
rect 29 447 45 481
rect 173 447 189 481
rect 29 400 189 447
rect 247 481 407 497
rect 247 447 263 481
rect 391 447 407 481
rect 247 400 407 447
rect 465 481 625 497
rect 465 447 481 481
rect 609 447 625 481
rect 465 400 625 447
rect 683 481 843 497
rect 683 447 699 481
rect 827 447 843 481
rect 683 400 843 447
rect 901 481 1061 497
rect 901 447 917 481
rect 1045 447 1061 481
rect 901 400 1061 447
rect 1119 481 1279 497
rect 1119 447 1135 481
rect 1263 447 1279 481
rect 1119 400 1279 447
rect -1279 -447 -1119 -400
rect -1279 -481 -1263 -447
rect -1135 -481 -1119 -447
rect -1279 -497 -1119 -481
rect -1061 -447 -901 -400
rect -1061 -481 -1045 -447
rect -917 -481 -901 -447
rect -1061 -497 -901 -481
rect -843 -447 -683 -400
rect -843 -481 -827 -447
rect -699 -481 -683 -447
rect -843 -497 -683 -481
rect -625 -447 -465 -400
rect -625 -481 -609 -447
rect -481 -481 -465 -447
rect -625 -497 -465 -481
rect -407 -447 -247 -400
rect -407 -481 -391 -447
rect -263 -481 -247 -447
rect -407 -497 -247 -481
rect -189 -447 -29 -400
rect -189 -481 -173 -447
rect -45 -481 -29 -447
rect -189 -497 -29 -481
rect 29 -447 189 -400
rect 29 -481 45 -447
rect 173 -481 189 -447
rect 29 -497 189 -481
rect 247 -447 407 -400
rect 247 -481 263 -447
rect 391 -481 407 -447
rect 247 -497 407 -481
rect 465 -447 625 -400
rect 465 -481 481 -447
rect 609 -481 625 -447
rect 465 -497 625 -481
rect 683 -447 843 -400
rect 683 -481 699 -447
rect 827 -481 843 -447
rect 683 -497 843 -481
rect 901 -447 1061 -400
rect 901 -481 917 -447
rect 1045 -481 1061 -447
rect 901 -497 1061 -481
rect 1119 -447 1279 -400
rect 1119 -481 1135 -447
rect 1263 -481 1279 -447
rect 1119 -497 1279 -481
<< polycont >>
rect -1263 447 -1135 481
rect -1045 447 -917 481
rect -827 447 -699 481
rect -609 447 -481 481
rect -391 447 -263 481
rect -173 447 -45 481
rect 45 447 173 481
rect 263 447 391 481
rect 481 447 609 481
rect 699 447 827 481
rect 917 447 1045 481
rect 1135 447 1263 481
rect -1263 -481 -1135 -447
rect -1045 -481 -917 -447
rect -827 -481 -699 -447
rect -609 -481 -481 -447
rect -391 -481 -263 -447
rect -173 -481 -45 -447
rect 45 -481 173 -447
rect 263 -481 391 -447
rect 481 -481 609 -447
rect 699 -481 827 -447
rect 917 -481 1045 -447
rect 1135 -481 1263 -447
<< locali >>
rect -1459 585 -1363 619
rect 1363 585 1459 619
rect -1459 523 -1425 585
rect 1425 523 1459 585
rect -1279 447 -1263 481
rect -1135 447 -1119 481
rect -1061 447 -1045 481
rect -917 447 -901 481
rect -843 447 -827 481
rect -699 447 -683 481
rect -625 447 -609 481
rect -481 447 -465 481
rect -407 447 -391 481
rect -263 447 -247 481
rect -189 447 -173 481
rect -45 447 -29 481
rect 29 447 45 481
rect 173 447 189 481
rect 247 447 263 481
rect 391 447 407 481
rect 465 447 481 481
rect 609 447 625 481
rect 683 447 699 481
rect 827 447 843 481
rect 901 447 917 481
rect 1045 447 1061 481
rect 1119 447 1135 481
rect 1263 447 1279 481
rect -1325 388 -1291 404
rect -1325 -404 -1291 -388
rect -1107 388 -1073 404
rect -1107 -404 -1073 -388
rect -889 388 -855 404
rect -889 -404 -855 -388
rect -671 388 -637 404
rect -671 -404 -637 -388
rect -453 388 -419 404
rect -453 -404 -419 -388
rect -235 388 -201 404
rect -235 -404 -201 -388
rect -17 388 17 404
rect -17 -404 17 -388
rect 201 388 235 404
rect 201 -404 235 -388
rect 419 388 453 404
rect 419 -404 453 -388
rect 637 388 671 404
rect 637 -404 671 -388
rect 855 388 889 404
rect 855 -404 889 -388
rect 1073 388 1107 404
rect 1073 -404 1107 -388
rect 1291 388 1325 404
rect 1291 -404 1325 -388
rect -1279 -481 -1263 -447
rect -1135 -481 -1119 -447
rect -1061 -481 -1045 -447
rect -917 -481 -901 -447
rect -843 -481 -827 -447
rect -699 -481 -683 -447
rect -625 -481 -609 -447
rect -481 -481 -465 -447
rect -407 -481 -391 -447
rect -263 -481 -247 -447
rect -189 -481 -173 -447
rect -45 -481 -29 -447
rect 29 -481 45 -447
rect 173 -481 189 -447
rect 247 -481 263 -447
rect 391 -481 407 -447
rect 465 -481 481 -447
rect 609 -481 625 -447
rect 683 -481 699 -447
rect 827 -481 843 -447
rect 901 -481 917 -447
rect 1045 -481 1061 -447
rect 1119 -481 1135 -447
rect 1263 -481 1279 -447
rect -1459 -585 -1425 -523
rect 1425 -585 1459 -523
rect -1459 -619 -1363 -585
rect 1363 -619 1459 -585
<< viali >>
rect -1263 447 -1135 481
rect -1045 447 -917 481
rect -827 447 -699 481
rect -609 447 -481 481
rect -391 447 -263 481
rect -173 447 -45 481
rect 45 447 173 481
rect 263 447 391 481
rect 481 447 609 481
rect 699 447 827 481
rect 917 447 1045 481
rect 1135 447 1263 481
rect -1325 -388 -1291 388
rect -1107 -388 -1073 388
rect -889 -388 -855 388
rect -671 -388 -637 388
rect -453 -388 -419 388
rect -235 -388 -201 388
rect -17 -388 17 388
rect 201 -388 235 388
rect 419 -388 453 388
rect 637 -388 671 388
rect 855 -388 889 388
rect 1073 -388 1107 388
rect 1291 -388 1325 388
rect -1263 -481 -1135 -447
rect -1045 -481 -917 -447
rect -827 -481 -699 -447
rect -609 -481 -481 -447
rect -391 -481 -263 -447
rect -173 -481 -45 -447
rect 45 -481 173 -447
rect 263 -481 391 -447
rect 481 -481 609 -447
rect 699 -481 827 -447
rect 917 -481 1045 -447
rect 1135 -481 1263 -447
<< metal1 >>
rect -1275 481 -1123 487
rect -1275 447 -1263 481
rect -1135 447 -1123 481
rect -1275 441 -1123 447
rect -1057 481 -905 487
rect -1057 447 -1045 481
rect -917 447 -905 481
rect -1057 441 -905 447
rect -839 481 -687 487
rect -839 447 -827 481
rect -699 447 -687 481
rect -839 441 -687 447
rect -621 481 -469 487
rect -621 447 -609 481
rect -481 447 -469 481
rect -621 441 -469 447
rect -403 481 -251 487
rect -403 447 -391 481
rect -263 447 -251 481
rect -403 441 -251 447
rect -185 481 -33 487
rect -185 447 -173 481
rect -45 447 -33 481
rect -185 441 -33 447
rect 33 481 185 487
rect 33 447 45 481
rect 173 447 185 481
rect 33 441 185 447
rect 251 481 403 487
rect 251 447 263 481
rect 391 447 403 481
rect 251 441 403 447
rect 469 481 621 487
rect 469 447 481 481
rect 609 447 621 481
rect 469 441 621 447
rect 687 481 839 487
rect 687 447 699 481
rect 827 447 839 481
rect 687 441 839 447
rect 905 481 1057 487
rect 905 447 917 481
rect 1045 447 1057 481
rect 905 441 1057 447
rect 1123 481 1275 487
rect 1123 447 1135 481
rect 1263 447 1275 481
rect 1123 441 1275 447
rect -1331 388 -1285 400
rect -1331 -388 -1325 388
rect -1291 -388 -1285 388
rect -1331 -400 -1285 -388
rect -1113 388 -1067 400
rect -1113 -388 -1107 388
rect -1073 -388 -1067 388
rect -1113 -400 -1067 -388
rect -895 388 -849 400
rect -895 -388 -889 388
rect -855 -388 -849 388
rect -895 -400 -849 -388
rect -677 388 -631 400
rect -677 -388 -671 388
rect -637 -388 -631 388
rect -677 -400 -631 -388
rect -459 388 -413 400
rect -459 -388 -453 388
rect -419 -388 -413 388
rect -459 -400 -413 -388
rect -241 388 -195 400
rect -241 -388 -235 388
rect -201 -388 -195 388
rect -241 -400 -195 -388
rect -23 388 23 400
rect -23 -388 -17 388
rect 17 -388 23 388
rect -23 -400 23 -388
rect 195 388 241 400
rect 195 -388 201 388
rect 235 -388 241 388
rect 195 -400 241 -388
rect 413 388 459 400
rect 413 -388 419 388
rect 453 -388 459 388
rect 413 -400 459 -388
rect 631 388 677 400
rect 631 -388 637 388
rect 671 -388 677 388
rect 631 -400 677 -388
rect 849 388 895 400
rect 849 -388 855 388
rect 889 -388 895 388
rect 849 -400 895 -388
rect 1067 388 1113 400
rect 1067 -388 1073 388
rect 1107 -388 1113 388
rect 1067 -400 1113 -388
rect 1285 388 1331 400
rect 1285 -388 1291 388
rect 1325 -388 1331 388
rect 1285 -400 1331 -388
rect -1275 -447 -1123 -441
rect -1275 -481 -1263 -447
rect -1135 -481 -1123 -447
rect -1275 -487 -1123 -481
rect -1057 -447 -905 -441
rect -1057 -481 -1045 -447
rect -917 -481 -905 -447
rect -1057 -487 -905 -481
rect -839 -447 -687 -441
rect -839 -481 -827 -447
rect -699 -481 -687 -447
rect -839 -487 -687 -481
rect -621 -447 -469 -441
rect -621 -481 -609 -447
rect -481 -481 -469 -447
rect -621 -487 -469 -481
rect -403 -447 -251 -441
rect -403 -481 -391 -447
rect -263 -481 -251 -447
rect -403 -487 -251 -481
rect -185 -447 -33 -441
rect -185 -481 -173 -447
rect -45 -481 -33 -447
rect -185 -487 -33 -481
rect 33 -447 185 -441
rect 33 -481 45 -447
rect 173 -481 185 -447
rect 33 -487 185 -481
rect 251 -447 403 -441
rect 251 -481 263 -447
rect 391 -481 403 -447
rect 251 -487 403 -481
rect 469 -447 621 -441
rect 469 -481 481 -447
rect 609 -481 621 -447
rect 469 -487 621 -481
rect 687 -447 839 -441
rect 687 -481 699 -447
rect 827 -481 839 -447
rect 687 -487 839 -481
rect 905 -447 1057 -441
rect 905 -481 917 -447
rect 1045 -481 1057 -447
rect 905 -487 1057 -481
rect 1123 -447 1275 -441
rect 1123 -481 1135 -447
rect 1263 -481 1275 -447
rect 1123 -487 1275 -481
<< properties >>
string FIXED_BBOX -1442 -602 1442 602
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 4 l 0.8 m 1 nf 12 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
