* Extracted by KLayout with SKY130 LVS runset on : 14/02/2025 00:58

.SUBCKT TOP
X$1 \$1 guard_ring_gen
X$2 \$1 vias_gen$1
X$3 \$2 \$1 \$1 \$1 pfet
X$4 \$1 \$1 \$2 \$1 pfet
X$5 \$1 \$1 \$2 \$1 pfet
X$6 \$2 \$1 \$1 \$1 pfet
X$7 \$2 \$2 \$1 \$1 pfet
X$8 \$1 \$1 \$18 \$2 \$2 \$1 pfet$1
X$9 \$2 \$2 \$1 \$1 pfet
X$10 \$1 \$1 \$18 \$2 \$2 \$1 pfet$1
X$11 \$1 \$2 \$2 \$1 pfet
X$12 \$1 \$2 \$2 \$1 pfet
X$13 \$2 vias_gen$3
X$14 \$2 vias_gen$3
X$15 \$2 vias_gen$3
X$16 \$2 vias_gen$3
X$17 \$2 vias_gen$5
X$18 \$2 vias_gen$5
X$19 \$2 vias_gen$5
X$20 \$2 vias_gen$5
X$21 \$2 vias_gen$5
X$22 \$2 vias_gen$5
X$23 \$2 vias_gen$5
X$24 \$2 vias_gen$5
X$25 \$2 vias_gen$5
X$26 \$2 vias_gen$5
X$27 \$2 vias_gen$5
X$28 \$2 vias_gen$5
X$29 \$2 vias_gen$5
X$30 \$2 vias_gen$5
X$31 \$2 vias_gen$5
X$32 \$2 vias_gen$5
M$1 \$1 \$1 \$2 \$1 sky130_fd_pr__pfet_g5v0d10v5 L=3 W=1.5 AS=0.45 AD=0.225
+ PS=3.6 PD=1.8
M$2 \$2 \$2 \$1 \$1 sky130_fd_pr__pfet_g5v0d10v5 L=3 W=1.5 AS=0.225 AD=0.225
+ PS=1.8 PD=1.8
M$3 \$1 \$2 \$18 \$1 sky130_fd_pr__pfet_g5v0d10v5 L=3 W=1.5 AS=0.225 AD=0.375
+ PS=1.8 PD=2
M$4 \$18 \$2 \$1 \$1 sky130_fd_pr__pfet_g5v0d10v5 L=3 W=1.5 AS=0.375 AD=0.225
+ PS=2 PD=1.8
M$5 \$1 \$2 \$2 \$1 sky130_fd_pr__pfet_g5v0d10v5 L=3 W=1.5 AS=0.225 AD=0.225
+ PS=1.8 PD=1.8
M$6 \$2 \$1 \$1 \$1 sky130_fd_pr__pfet_g5v0d10v5 L=3 W=1.5 AS=0.225 AD=0.45
+ PS=1.8 PD=3.6
M$7 \$1 \$1 \$2 \$1 sky130_fd_pr__pfet_g5v0d10v5 L=3 W=1.5 AS=0.45 AD=0.225
+ PS=3.6 PD=1.8
M$8 \$2 \$2 \$1 \$1 sky130_fd_pr__pfet_g5v0d10v5 L=3 W=1.5 AS=0.225 AD=0.225
+ PS=1.8 PD=1.8
M$9 \$1 \$2 \$18 \$1 sky130_fd_pr__pfet_g5v0d10v5 L=3 W=1.5 AS=0.225 AD=0.375
+ PS=1.8 PD=2
M$10 \$18 \$2 \$1 \$1 sky130_fd_pr__pfet_g5v0d10v5 L=3 W=1.5 AS=0.375 AD=0.225
+ PS=2 PD=1.8
M$11 \$1 \$2 \$2 \$1 sky130_fd_pr__pfet_g5v0d10v5 L=3 W=1.5 AS=0.225 AD=0.225
+ PS=1.8 PD=1.8
M$12 \$2 \$1 \$1 \$1 sky130_fd_pr__pfet_g5v0d10v5 L=3 W=1.5 AS=0.225 AD=0.45
+ PS=1.8 PD=3.6
.ENDS TOP

.SUBCKT vias_gen$5 \$1
.ENDS vias_gen$5

.SUBCKT vias_gen$3 \$1
.ENDS vias_gen$3

.SUBCKT vias_gen$1 \$1
.ENDS vias_gen$1

.SUBCKT guard_ring_gen \$2
.ENDS guard_ring_gen

.SUBCKT pfet$1 \$1 \$2 \$3 \$4 \$5 \$6
.ENDS pfet$1

.SUBCKT pfet \$1 \$2 \$3 \$4
.ENDS pfet
