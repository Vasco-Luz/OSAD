** sch_path: /foss/designs/OSAD/Learning/single_ended_amplifiers/Design_and_Analysis_of_Two-Stage_CMOS_Operational_Amplifier_for_Fluorescence_Signal_Processing_ihp130_3_3V/transcondutance/design.sch
**.subckt design
V1 VDD GND 3.3
V2 VSS GND 0
XM2 VB1 VB1 VDD VDD sg13_hv_pmos w=1.0u l=2u ng=2 m=2
XM1 VB2 VB1 VDD VDD sg13_hv_pmos w=1.0u l=2u ng=2 m=2
XM3 VB1 VB2 net3 VSS sg13_hv_nmos w=1.0u l=2u ng=2 m=2
XM4 VB2 VB2 net1 VSS sg13_hv_nmos w=1.0u l=2u ng=2 m=2
XM5 net4 net1 net2 VSS sg13_hv_nmos w=2u l=2u ng=2 m=8
XM6 net1 net1 VSS VSS sg13_hv_nmos w=2u l=2u ng=2 m=2
Vmeas net3 net4 0
.save i(vmeas)
XR1 VSS net2 rhigh w=0.5e-6 l=5.9e-6 m=1 b=0
XM7 net5 VB1 VDD VDD sg13_hv_pmos w=1.0u l=2u ng=2 m=2
Vmeas1 net5 net6 0
.save i(vmeas1)
V3 net6 GND 3.3
**** begin user architecture code

.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerRES.lib res_typ_stat



.param mm_ok=1
.param mc_ok=1
.param temp=27
.control
save all
dc temp -50 125 1
plot i(Vmeas)
dc V3 0 3.3 0.001
plot i(Vmeas1)


.endc



.lib cornerMOShv.lib mos_tt_stat

**** end user architecture code
**.ends
.GLOBAL GND
.end
