magic
tech sky130A
magscale 1 2
timestamp 1740356695
<< error_p >>
rect -1403 -131 -1345 69
rect -945 -131 -887 69
rect -487 -131 -429 69
rect -29 -131 29 69
rect 429 -131 487 69
rect 887 -131 945 69
rect 1345 -131 1403 69
rect 1803 -131 1861 69
rect 2261 -131 2319 69
<< mvnmos >>
rect -2261 -131 -1861 69
rect -1803 -131 -1403 69
rect -1345 -131 -945 69
rect -887 -131 -487 69
rect -429 -131 -29 69
rect 29 -131 429 69
rect 487 -131 887 69
rect 945 -131 1345 69
rect 1403 -131 1803 69
rect 1861 -131 2261 69
<< mvndiff >>
rect -2319 57 -2261 69
rect -2319 -119 -2307 57
rect -2273 -119 -2261 57
rect -2319 -131 -2261 -119
rect -1861 57 -1803 69
rect -1861 -119 -1849 57
rect -1815 -119 -1803 57
rect -1861 -131 -1803 -119
rect -1403 57 -1345 69
rect -1403 -119 -1391 57
rect -1357 -119 -1345 57
rect -1403 -131 -1345 -119
rect -945 57 -887 69
rect -945 -119 -933 57
rect -899 -119 -887 57
rect -945 -131 -887 -119
rect -487 57 -429 69
rect -487 -119 -475 57
rect -441 -119 -429 57
rect -487 -131 -429 -119
rect -29 57 29 69
rect -29 -119 -17 57
rect 17 -119 29 57
rect -29 -131 29 -119
rect 429 57 487 69
rect 429 -119 441 57
rect 475 -119 487 57
rect 429 -131 487 -119
rect 887 57 945 69
rect 887 -119 899 57
rect 933 -119 945 57
rect 887 -131 945 -119
rect 1345 57 1403 69
rect 1345 -119 1357 57
rect 1391 -119 1403 57
rect 1345 -131 1403 -119
rect 1803 57 1861 69
rect 1803 -119 1815 57
rect 1849 -119 1861 57
rect 1803 -131 1861 -119
rect 2261 57 2319 69
rect 2261 -119 2273 57
rect 2307 -119 2319 57
rect 2261 -131 2319 -119
<< mvndiffc >>
rect -2307 -119 -2273 57
rect -1849 -119 -1815 57
rect -1391 -119 -1357 57
rect -933 -119 -899 57
rect -475 -119 -441 57
rect -17 -119 17 57
rect 441 -119 475 57
rect 899 -119 933 57
rect 1357 -119 1391 57
rect 1815 -119 1849 57
rect 2273 -119 2307 57
<< poly >>
rect -2224 141 -1898 157
rect -2224 124 -2208 141
rect -2261 107 -2208 124
rect -1914 124 -1898 141
rect -1766 141 -1440 157
rect -1766 124 -1750 141
rect -1914 107 -1861 124
rect -2261 69 -1861 107
rect -1803 107 -1750 124
rect -1456 124 -1440 141
rect -1308 141 -982 157
rect -1308 124 -1292 141
rect -1456 107 -1403 124
rect -1803 69 -1403 107
rect -1345 107 -1292 124
rect -998 124 -982 141
rect -850 141 -524 157
rect -850 124 -834 141
rect -998 107 -945 124
rect -1345 69 -945 107
rect -887 107 -834 124
rect -540 124 -524 141
rect -392 141 -66 157
rect -392 124 -376 141
rect -540 107 -487 124
rect -887 69 -487 107
rect -429 107 -376 124
rect -82 124 -66 141
rect 66 141 392 157
rect 66 124 82 141
rect -82 107 -29 124
rect -429 69 -29 107
rect 29 107 82 124
rect 376 124 392 141
rect 524 141 850 157
rect 524 124 540 141
rect 376 107 429 124
rect 29 69 429 107
rect 487 107 540 124
rect 834 124 850 141
rect 982 141 1308 157
rect 982 124 998 141
rect 834 107 887 124
rect 487 69 887 107
rect 945 107 998 124
rect 1292 124 1308 141
rect 1440 141 1766 157
rect 1440 124 1456 141
rect 1292 107 1345 124
rect 945 69 1345 107
rect 1403 107 1456 124
rect 1750 124 1766 141
rect 1898 141 2224 157
rect 1898 124 1914 141
rect 1750 107 1803 124
rect 1403 69 1803 107
rect 1861 107 1914 124
rect 2208 124 2224 141
rect 2208 107 2261 124
rect 1861 69 2261 107
rect -2261 -157 -1861 -131
rect -1803 -157 -1403 -131
rect -1345 -157 -945 -131
rect -887 -157 -487 -131
rect -429 -157 -29 -131
rect 29 -157 429 -131
rect 487 -157 887 -131
rect 945 -157 1345 -131
rect 1403 -157 1803 -131
rect 1861 -157 2261 -131
<< polycont >>
rect -2208 107 -1914 141
rect -1750 107 -1456 141
rect -1292 107 -998 141
rect -834 107 -540 141
rect -376 107 -82 141
rect 82 107 376 141
rect 540 107 834 141
rect 998 107 1292 141
rect 1456 107 1750 141
rect 1914 107 2208 141
<< locali >>
rect -2224 107 -2208 141
rect -1914 107 -1898 141
rect -1766 107 -1750 141
rect -1456 107 -1440 141
rect -1308 107 -1292 141
rect -998 107 -982 141
rect -850 107 -834 141
rect -540 107 -524 141
rect -392 107 -376 141
rect -82 107 -66 141
rect 66 107 82 141
rect 376 107 392 141
rect 524 107 540 141
rect 834 107 850 141
rect 982 107 998 141
rect 1292 107 1308 141
rect 1440 107 1456 141
rect 1750 107 1766 141
rect 1898 107 1914 141
rect 2208 107 2224 141
rect -2307 57 -2273 73
rect -2307 -135 -2273 -119
rect -1849 57 -1815 73
rect -1849 -135 -1815 -119
rect -1391 57 -1357 73
rect -1391 -135 -1357 -119
rect -933 57 -899 73
rect -933 -135 -899 -119
rect -475 57 -441 73
rect -475 -135 -441 -119
rect -17 57 17 73
rect -17 -135 17 -119
rect 441 57 475 73
rect 441 -135 475 -119
rect 899 57 933 73
rect 899 -135 933 -119
rect 1357 57 1391 73
rect 1357 -135 1391 -119
rect 1815 57 1849 73
rect 1815 -135 1849 -119
rect 2273 57 2307 73
rect 2273 -135 2307 -119
<< viali >>
rect -2208 107 -1914 141
rect -1750 107 -1456 141
rect -1292 107 -998 141
rect -834 107 -540 141
rect -376 107 -82 141
rect 82 107 376 141
rect 540 107 834 141
rect 998 107 1292 141
rect 1456 107 1750 141
rect 1914 107 2208 141
rect -2307 -119 -2273 57
rect -1849 -119 -1815 57
rect -1391 -119 -1357 57
rect -933 -119 -899 57
rect -475 -119 -441 57
rect -17 -119 17 57
rect 441 -119 475 57
rect 899 -119 933 57
rect 1357 -119 1391 57
rect 1815 -119 1849 57
rect 2273 -119 2307 57
<< metal1 >>
rect -2220 141 -1902 147
rect -2220 107 -2208 141
rect -1914 107 -1902 141
rect -2220 101 -1902 107
rect -1762 141 -1444 147
rect -1762 107 -1750 141
rect -1456 107 -1444 141
rect -1762 101 -1444 107
rect -1304 141 -986 147
rect -1304 107 -1292 141
rect -998 107 -986 141
rect -1304 101 -986 107
rect -846 141 -528 147
rect -846 107 -834 141
rect -540 107 -528 141
rect -846 101 -528 107
rect -388 141 -70 147
rect -388 107 -376 141
rect -82 107 -70 141
rect -388 101 -70 107
rect 70 141 388 147
rect 70 107 82 141
rect 376 107 388 141
rect 70 101 388 107
rect 528 141 846 147
rect 528 107 540 141
rect 834 107 846 141
rect 528 101 846 107
rect 986 141 1304 147
rect 986 107 998 141
rect 1292 107 1304 141
rect 986 101 1304 107
rect 1444 141 1762 147
rect 1444 107 1456 141
rect 1750 107 1762 141
rect 1444 101 1762 107
rect 1902 141 2220 147
rect 1902 107 1914 141
rect 2208 107 2220 141
rect 1902 101 2220 107
rect -2313 57 -2267 69
rect -2313 -119 -2307 57
rect -2273 -119 -2267 57
rect -2313 -131 -2267 -119
rect -1855 57 -1809 69
rect -1855 -119 -1849 57
rect -1815 -119 -1809 57
rect -1855 -131 -1809 -119
rect -1397 57 -1351 69
rect -1397 -119 -1391 57
rect -1357 -119 -1351 57
rect -1397 -131 -1351 -119
rect -939 57 -893 69
rect -939 -119 -933 57
rect -899 -119 -893 57
rect -939 -131 -893 -119
rect -481 57 -435 69
rect -481 -119 -475 57
rect -441 -119 -435 57
rect -481 -131 -435 -119
rect -23 57 23 69
rect -23 -119 -17 57
rect 17 -119 23 57
rect -23 -131 23 -119
rect 435 57 481 69
rect 435 -119 441 57
rect 475 -119 481 57
rect 435 -131 481 -119
rect 893 57 939 69
rect 893 -119 899 57
rect 933 -119 939 57
rect 893 -131 939 -119
rect 1351 57 1397 69
rect 1351 -119 1357 57
rect 1391 -119 1397 57
rect 1351 -131 1397 -119
rect 1809 57 1855 69
rect 1809 -119 1815 57
rect 1849 -119 1855 57
rect 1809 -131 1855 -119
rect 2267 57 2313 69
rect 2267 -119 2273 57
rect 2307 -119 2313 57
rect 2267 -131 2313 -119
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 1 l 2 m 1 nf 10 diffcov 100 polycov 80 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 80 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 80 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
