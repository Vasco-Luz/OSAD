magic
tech sky130A
magscale 1 2
timestamp 1693699723
<< nwell >>
rect -1537 -662 1537 662
<< mvpmos >>
rect -1279 -436 -1119 364
rect -1061 -436 -901 364
rect -843 -436 -683 364
rect -625 -436 -465 364
rect -407 -436 -247 364
rect -189 -436 -29 364
rect 29 -436 189 364
rect 247 -436 407 364
rect 465 -436 625 364
rect 683 -436 843 364
rect 901 -436 1061 364
rect 1119 -436 1279 364
<< mvpdiff >>
rect -1337 352 -1279 364
rect -1337 -424 -1325 352
rect -1291 -424 -1279 352
rect -1337 -436 -1279 -424
rect -1119 352 -1061 364
rect -1119 -424 -1107 352
rect -1073 -424 -1061 352
rect -1119 -436 -1061 -424
rect -901 352 -843 364
rect -901 -424 -889 352
rect -855 -424 -843 352
rect -901 -436 -843 -424
rect -683 352 -625 364
rect -683 -424 -671 352
rect -637 -424 -625 352
rect -683 -436 -625 -424
rect -465 352 -407 364
rect -465 -424 -453 352
rect -419 -424 -407 352
rect -465 -436 -407 -424
rect -247 352 -189 364
rect -247 -424 -235 352
rect -201 -424 -189 352
rect -247 -436 -189 -424
rect -29 352 29 364
rect -29 -424 -17 352
rect 17 -424 29 352
rect -29 -436 29 -424
rect 189 352 247 364
rect 189 -424 201 352
rect 235 -424 247 352
rect 189 -436 247 -424
rect 407 352 465 364
rect 407 -424 419 352
rect 453 -424 465 352
rect 407 -436 465 -424
rect 625 352 683 364
rect 625 -424 637 352
rect 671 -424 683 352
rect 625 -436 683 -424
rect 843 352 901 364
rect 843 -424 855 352
rect 889 -424 901 352
rect 843 -436 901 -424
rect 1061 352 1119 364
rect 1061 -424 1073 352
rect 1107 -424 1119 352
rect 1061 -436 1119 -424
rect 1279 352 1337 364
rect 1279 -424 1291 352
rect 1325 -424 1337 352
rect 1279 -436 1337 -424
<< mvpdiffc >>
rect -1325 -424 -1291 352
rect -1107 -424 -1073 352
rect -889 -424 -855 352
rect -671 -424 -637 352
rect -453 -424 -419 352
rect -235 -424 -201 352
rect -17 -424 17 352
rect 201 -424 235 352
rect 419 -424 453 352
rect 637 -424 671 352
rect 855 -424 889 352
rect 1073 -424 1107 352
rect 1291 -424 1325 352
<< mvnsubdiff >>
rect -1471 584 1471 596
rect -1471 550 -1363 584
rect 1363 550 1471 584
rect -1471 538 1471 550
rect -1471 488 -1413 538
rect -1471 -488 -1459 488
rect -1425 -488 -1413 488
rect 1413 488 1471 538
rect -1471 -538 -1413 -488
rect 1413 -488 1425 488
rect 1459 -488 1471 488
rect 1413 -538 1471 -488
rect -1471 -550 1471 -538
rect -1471 -584 -1363 -550
rect 1363 -584 1471 -550
rect -1471 -596 1471 -584
<< mvnsubdiffcont >>
rect -1363 550 1363 584
rect -1459 -488 -1425 488
rect 1425 -488 1459 488
rect -1363 -584 1363 -550
<< poly >>
rect -1260 445 -1138 461
rect -1260 428 -1244 445
rect -1279 411 -1244 428
rect -1154 428 -1138 445
rect -1042 445 -920 461
rect -1042 428 -1026 445
rect -1154 411 -1119 428
rect -1279 364 -1119 411
rect -1061 411 -1026 428
rect -936 428 -920 445
rect -824 445 -702 461
rect -824 428 -808 445
rect -936 411 -901 428
rect -1061 364 -901 411
rect -843 411 -808 428
rect -718 428 -702 445
rect -606 445 -484 461
rect -606 428 -590 445
rect -718 411 -683 428
rect -843 364 -683 411
rect -625 411 -590 428
rect -500 428 -484 445
rect -388 445 -266 461
rect -388 428 -372 445
rect -500 411 -465 428
rect -625 364 -465 411
rect -407 411 -372 428
rect -282 428 -266 445
rect -170 445 -48 461
rect -170 428 -154 445
rect -282 411 -247 428
rect -407 364 -247 411
rect -189 411 -154 428
rect -64 428 -48 445
rect 48 445 170 461
rect 48 428 64 445
rect -64 411 -29 428
rect -189 364 -29 411
rect 29 411 64 428
rect 154 428 170 445
rect 266 445 388 461
rect 266 428 282 445
rect 154 411 189 428
rect 29 364 189 411
rect 247 411 282 428
rect 372 428 388 445
rect 484 445 606 461
rect 484 428 500 445
rect 372 411 407 428
rect 247 364 407 411
rect 465 411 500 428
rect 590 428 606 445
rect 702 445 824 461
rect 702 428 718 445
rect 590 411 625 428
rect 465 364 625 411
rect 683 411 718 428
rect 808 428 824 445
rect 920 445 1042 461
rect 920 428 936 445
rect 808 411 843 428
rect 683 364 843 411
rect 901 411 936 428
rect 1026 428 1042 445
rect 1138 445 1260 461
rect 1138 428 1154 445
rect 1026 411 1061 428
rect 901 364 1061 411
rect 1119 411 1154 428
rect 1244 428 1260 445
rect 1244 411 1279 428
rect 1119 364 1279 411
rect -1279 -462 -1119 -436
rect -1061 -462 -901 -436
rect -843 -462 -683 -436
rect -625 -462 -465 -436
rect -407 -462 -247 -436
rect -189 -462 -29 -436
rect 29 -462 189 -436
rect 247 -462 407 -436
rect 465 -462 625 -436
rect 683 -462 843 -436
rect 901 -462 1061 -436
rect 1119 -462 1279 -436
<< polycont >>
rect -1244 411 -1154 445
rect -1026 411 -936 445
rect -808 411 -718 445
rect -590 411 -500 445
rect -372 411 -282 445
rect -154 411 -64 445
rect 64 411 154 445
rect 282 411 372 445
rect 500 411 590 445
rect 718 411 808 445
rect 936 411 1026 445
rect 1154 411 1244 445
<< locali >>
rect -1459 550 -1363 584
rect 1363 550 1459 584
rect -1459 488 -1425 550
rect 1425 488 1459 550
rect -1260 411 -1244 445
rect -1154 411 -1138 445
rect -1042 411 -1026 445
rect -936 411 -920 445
rect -824 411 -808 445
rect -718 411 -702 445
rect -606 411 -590 445
rect -500 411 -484 445
rect -388 411 -372 445
rect -282 411 -266 445
rect -170 411 -154 445
rect -64 411 -48 445
rect 48 411 64 445
rect 154 411 170 445
rect 266 411 282 445
rect 372 411 388 445
rect 484 411 500 445
rect 590 411 606 445
rect 702 411 718 445
rect 808 411 824 445
rect 920 411 936 445
rect 1026 411 1042 445
rect 1138 411 1154 445
rect 1244 411 1260 445
rect -1325 352 -1291 368
rect -1325 -440 -1291 -424
rect -1107 352 -1073 368
rect -1107 -440 -1073 -424
rect -889 352 -855 368
rect -889 -440 -855 -424
rect -671 352 -637 368
rect -671 -440 -637 -424
rect -453 352 -419 368
rect -453 -440 -419 -424
rect -235 352 -201 368
rect -235 -440 -201 -424
rect -17 352 17 368
rect -17 -440 17 -424
rect 201 352 235 368
rect 201 -440 235 -424
rect 419 352 453 368
rect 419 -440 453 -424
rect 637 352 671 368
rect 637 -440 671 -424
rect 855 352 889 368
rect 855 -440 889 -424
rect 1073 352 1107 368
rect 1073 -440 1107 -424
rect 1291 352 1325 368
rect 1291 -440 1325 -424
rect -1459 -550 -1425 -488
rect 1425 -550 1459 -488
rect -1459 -584 -1363 -550
rect 1363 -584 1459 -550
<< viali >>
rect -1244 411 -1154 445
rect -1026 411 -936 445
rect -808 411 -718 445
rect -590 411 -500 445
rect -372 411 -282 445
rect -154 411 -64 445
rect 64 411 154 445
rect 282 411 372 445
rect 500 411 590 445
rect 718 411 808 445
rect 936 411 1026 445
rect 1154 411 1244 445
rect -1325 -424 -1291 352
rect -1107 -424 -1073 352
rect -889 -424 -855 352
rect -671 -424 -637 352
rect -453 -424 -419 352
rect -235 -424 -201 352
rect -17 -424 17 352
rect 201 -424 235 352
rect 419 -424 453 352
rect 637 -424 671 352
rect 855 -424 889 352
rect 1073 -424 1107 352
rect 1291 -424 1325 352
<< metal1 >>
rect -1256 445 -1142 451
rect -1256 411 -1244 445
rect -1154 411 -1142 445
rect -1256 405 -1142 411
rect -1038 445 -924 451
rect -1038 411 -1026 445
rect -936 411 -924 445
rect -1038 405 -924 411
rect -820 445 -706 451
rect -820 411 -808 445
rect -718 411 -706 445
rect -820 405 -706 411
rect -602 445 -488 451
rect -602 411 -590 445
rect -500 411 -488 445
rect -602 405 -488 411
rect -384 445 -270 451
rect -384 411 -372 445
rect -282 411 -270 445
rect -384 405 -270 411
rect -166 445 -52 451
rect -166 411 -154 445
rect -64 411 -52 445
rect -166 405 -52 411
rect 52 445 166 451
rect 52 411 64 445
rect 154 411 166 445
rect 52 405 166 411
rect 270 445 384 451
rect 270 411 282 445
rect 372 411 384 445
rect 270 405 384 411
rect 488 445 602 451
rect 488 411 500 445
rect 590 411 602 445
rect 488 405 602 411
rect 706 445 820 451
rect 706 411 718 445
rect 808 411 820 445
rect 706 405 820 411
rect 924 445 1038 451
rect 924 411 936 445
rect 1026 411 1038 445
rect 924 405 1038 411
rect 1142 445 1256 451
rect 1142 411 1154 445
rect 1244 411 1256 445
rect 1142 405 1256 411
rect -1331 352 -1285 364
rect -1331 -424 -1325 352
rect -1291 -424 -1285 352
rect -1331 -436 -1285 -424
rect -1113 352 -1067 364
rect -1113 -424 -1107 352
rect -1073 -424 -1067 352
rect -1113 -436 -1067 -424
rect -895 352 -849 364
rect -895 -424 -889 352
rect -855 -424 -849 352
rect -895 -436 -849 -424
rect -677 352 -631 364
rect -677 -424 -671 352
rect -637 -424 -631 352
rect -677 -436 -631 -424
rect -459 352 -413 364
rect -459 -424 -453 352
rect -419 -424 -413 352
rect -459 -436 -413 -424
rect -241 352 -195 364
rect -241 -424 -235 352
rect -201 -424 -195 352
rect -241 -436 -195 -424
rect -23 352 23 364
rect -23 -424 -17 352
rect 17 -424 23 352
rect -23 -436 23 -424
rect 195 352 241 364
rect 195 -424 201 352
rect 235 -424 241 352
rect 195 -436 241 -424
rect 413 352 459 364
rect 413 -424 419 352
rect 453 -424 459 352
rect 413 -436 459 -424
rect 631 352 677 364
rect 631 -424 637 352
rect 671 -424 677 352
rect 631 -436 677 -424
rect 849 352 895 364
rect 849 -424 855 352
rect 889 -424 895 352
rect 849 -436 895 -424
rect 1067 352 1113 364
rect 1067 -424 1073 352
rect 1107 -424 1113 352
rect 1067 -436 1113 -424
rect 1285 352 1331 364
rect 1285 -424 1291 352
rect 1325 -424 1331 352
rect 1285 -436 1331 -424
<< properties >>
string FIXED_BBOX -1442 -567 1442 567
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 4 l 0.8 m 1 nf 12 diffcov 100 polycov 70 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 70 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
