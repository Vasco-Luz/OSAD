* Extracted by KLayout with SKY130 LVS runset on : 04/03/2025 01:44

.SUBCKT upper_nmos_current_mirror VSS
M$1 \$3 \$3 \$1 VSS sky130_fd_pr__nfet_g5v0d10v5 L=2000000 W=4000000 AS=1.1e+12
+ AD=1.1e+12 PS=8200000 PD=8200000
M$2 \$1 \$1 \$9 VSS sky130_fd_pr__nfet_g5v0d10v5 L=2000000 W=4000000 AS=1e+12
+ AD=1e+12 PS=6000000 PD=6000000
M$3 \$9 \$3 \$3 VSS sky130_fd_pr__nfet_g5v0d10v5 L=2000000 W=4000000 AS=1e+12
+ AD=1e+12 PS=6000000 PD=6000000
M$4 \$3 \$3 \$17 VSS sky130_fd_pr__nfet_g5v0d10v5 L=2000000 W=4000000 AS=1e+12
+ AD=1e+12 PS=6000000 PD=6000000
M$5 \$17 \$1 \$11 VSS sky130_fd_pr__nfet_g5v0d10v5 L=2000000 W=4000000 AS=1e+12
+ AD=1e+12 PS=6000000 PD=6000000
.ENDS upper_nmos_current_mirror
