** sch_path: /foss/designs/OSAD/Learning/single_ended_amplifiers/Design_and_Analysis_of_Two-Stage_CMOS_Operational_Amplifier_for_Fluorescence_Signal_Processing_sky130_5V/klayout_layout/upper_nmos_current_mirror.sch
.subckt upper_nmos_current_mirror VSS IA IB IC ID
*.PININFO VSS:B IA:B IB:B IC:B ID:B
M9 IA IB IC VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W='1 * 2 ' nf=2 m=2
M10 IB IB ID VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W='1 * 2 ' nf=2 m=2
M1 IA VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W='1 * 1 ' nf=1 m=4
M2 IB VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W='1 * 1 ' nf=1 m=4
M3 ID VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W='1 * 1 ' nf=1 m=4
.ends
.end
