** sch_path: /home/vasco/PDK/ihp-sg13g2/libs.tech/xschem/sg13g2_tests/dc_ntap1.sch
**.subckt dc_ntap1
Vres Vcc GND 1.5
XR1 GND net1 ntap1
Vmeas Vcc net1 0
.save i(vmeas)
**** begin user architecture code

.lib /home/vasco/PDK/ihp-sg13g2/libs.tech/ngspice/models/cornerRES.lib res_typ



.param temp=27
.control
save all
op
print Vcc/I(Vr)
reset
dc Vres 0 3 0.01
write dc_ntap1.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
