magic
tech sky130A
magscale 1 2
timestamp 1693784648
<< nwell >>
rect -428 -657 428 657
<< nsubdiff >>
rect -392 587 -296 621
rect 296 587 392 621
rect -392 525 -358 587
rect 358 525 392 587
rect -392 -587 -358 -525
rect 358 -587 392 -525
rect -392 -621 -296 -587
rect 296 -621 392 -587
<< nsubdiffcont >>
rect -296 587 296 621
rect -392 -525 -358 525
rect 358 -525 392 525
rect -296 -621 296 -587
<< xpolycontact >>
rect -201 50 -131 482
rect -201 -482 -131 -50
rect -35 50 35 482
rect -35 -482 35 -50
rect 131 50 201 482
rect 131 -482 201 -50
<< ppolyres >>
rect -201 -50 -131 50
rect -35 -50 35 50
rect 131 -50 201 50
<< locali >>
rect -392 587 -296 621
rect 296 587 392 621
rect -392 525 -358 587
rect 358 525 392 587
rect -392 -587 -358 -525
rect 358 -587 392 -525
rect -392 -621 -296 -587
rect 296 -621 392 -587
<< viali >>
rect -185 67 -147 464
rect -19 67 19 464
rect 147 67 185 464
rect -185 -464 -147 -67
rect -19 -464 19 -67
rect 147 -464 185 -67
<< metal1 >>
rect -191 464 -141 476
rect -191 67 -185 464
rect -147 67 -141 464
rect -191 55 -141 67
rect -25 464 25 476
rect -25 67 -19 464
rect 19 67 25 464
rect -25 55 25 67
rect 141 464 191 476
rect 141 67 147 464
rect 185 67 191 464
rect 141 55 191 67
rect -191 -67 -141 -55
rect -191 -464 -185 -67
rect -147 -464 -141 -67
rect -191 -476 -141 -464
rect -25 -67 25 -55
rect -25 -464 -19 -67
rect 19 -464 25 -67
rect -25 -476 25 -464
rect 141 -67 191 -55
rect 141 -464 147 -67
rect 185 -464 191 -67
rect 141 -476 191 -464
<< properties >>
string FIXED_BBOX -375 -604 375 604
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.35 l 0.5 m 1 nx 3 wmin 0.350 lmin 0.50 rho 319.8 val 1.57k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 1 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
