magic
tech sky130A
magscale 1 2
timestamp 1740491809
<< mvpsubdiff >>
rect -2491 1967 -2431 2001
rect 2167 1967 2227 2001
rect -2491 1941 -2457 1967
rect -2491 -2151 -2457 -2125
rect 2193 1941 2227 1967
rect 2193 -2151 2227 -2125
rect -2491 -2185 -2431 -2151
rect 2167 -2185 2227 -2151
<< mvpsubdiffcont >>
rect -2431 1967 2167 2001
rect -2491 -2125 -2457 1941
rect 2193 -2125 2227 1941
rect -2431 -2185 2167 -2151
<< locali >>
rect -2862 2001 -2456 2008
rect -2862 1967 -2431 2001
rect 2167 1967 2227 2001
rect -2862 1941 -2456 1967
rect -2862 -2125 -2491 1941
rect -2457 -2125 -2456 1941
rect -2862 -2151 -2456 -2125
rect 2193 1941 2227 1967
rect 2193 -2151 2227 -2125
rect -2862 -2176 -2431 -2151
rect -2491 -2185 -2431 -2176
rect 2167 -2185 2227 -2151
<< metal3 >>
rect -334 2268 -234 2284
rect 1878 2268 1978 2282
rect -334 2204 -316 2268
rect -252 2266 1978 2268
rect -252 2204 1896 2266
rect -334 2184 -234 2204
rect 1878 2202 1896 2204
rect 1960 2202 1978 2266
rect 1878 2184 1978 2202
rect -1414 2124 -1314 2140
rect -1414 2060 -1396 2124
rect -1332 2108 898 2124
rect -1332 2060 816 2108
rect -1414 2040 -1314 2060
rect 798 2044 816 2060
rect 880 2044 898 2108
rect 798 2024 898 2044
<< via3 >>
rect -316 2204 -252 2268
rect 1896 2202 1960 2266
rect -1396 2060 -1332 2124
rect 816 2044 880 2108
<< metal4 >>
rect -338 2268 -234 2284
rect -338 2204 -316 2268
rect -252 2204 -234 2268
rect -1418 2124 -1314 2140
rect -1418 2060 -1396 2124
rect -1332 2060 -1314 2124
rect -1418 1786 -1314 2060
rect -338 1808 -234 2204
rect 1874 2266 1978 2282
rect 1874 2202 1896 2266
rect 1960 2202 1978 2266
rect 794 2108 898 2124
rect 794 2044 816 2108
rect 880 2044 898 2108
rect 794 1778 898 2044
rect 1874 1830 1978 2202
use sky130_fd_pr__cap_mim_m3_1_7PSTXW  sky130_fd_pr__cap_mim_m3_1_7PSTXW_0
timestamp 1740488682
transform 1 0 -114 0 1 -46
box -2092 -1920 2092 1920
<< labels >>
flabel locali -2736 -734 -2656 -636 0 FreeSans 1600 0 0 0 VSS
port 1 nsew
flabel metal3 -896 2084 -854 2096 0 FreeSans 1600 0 0 0 Ib
port 3 nsew
flabel metal3 506 2234 558 2250 0 FreeSans 1600 0 0 0 VOUT
port 5 nsew
<< end >>
