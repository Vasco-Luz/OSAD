magic
tech sky130A
magscale 1 2
timestamp 1740484998
<< mvnmos >>
rect -100 -431 100 369
<< mvndiff >>
rect -158 357 -100 369
rect -158 -419 -146 357
rect -112 -419 -100 357
rect -158 -431 -100 -419
rect 100 357 158 369
rect 100 -419 112 357
rect 146 -419 158 357
rect 100 -431 158 -419
<< mvndiffc >>
rect -146 -419 -112 357
rect 112 -419 146 357
<< poly >>
rect -83 441 83 457
rect -83 424 -67 441
rect -100 407 -67 424
rect 67 424 83 441
rect 67 407 100 424
rect -100 369 100 407
rect -100 -457 100 -431
<< polycont >>
rect -67 407 67 441
<< locali >>
rect -83 407 -67 441
rect 67 407 83 441
rect -146 357 -112 373
rect -146 -435 -112 -419
rect 112 357 146 373
rect 112 -435 146 -419
<< viali >>
rect -67 407 67 441
rect -146 -419 -112 357
rect 112 -419 146 357
<< metal1 >>
rect -79 441 79 447
rect -79 407 -67 441
rect 67 407 79 441
rect -79 401 79 407
rect -152 357 -106 369
rect -152 -419 -146 357
rect -112 -419 -106 357
rect -152 -431 -106 -419
rect 106 357 152 369
rect 106 -419 112 357
rect 146 -419 152 357
rect 106 -431 152 -419
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4 l 1 m 1 nf 1 diffcov 100 polycov 80 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 80 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
