magic
tech sky130A
magscale 1 2
timestamp 1738973162
<< nwell >>
rect -841 -155 2273 1093
<< mvnsubdiff >>
rect -775 993 -715 1027
rect 2147 993 2207 1027
rect -775 967 -741 993
rect -775 -55 -741 -29
rect 2173 967 2207 993
rect 2173 -55 2207 -29
rect -775 -89 -715 -55
rect 2147 -89 2207 -55
<< mvnsubdiffcont >>
rect -715 993 2147 1027
rect -775 -29 -741 967
rect 2173 -29 2207 967
rect -715 -89 2147 -55
<< locali >>
rect -775 994 -746 1027
rect -775 993 -715 994
rect 2147 993 2207 1027
rect -775 967 -741 993
rect -775 -55 -741 -29
rect 2173 967 2207 993
rect 2173 -55 2207 -29
rect -775 -89 -715 -55
rect 2147 -89 2207 -55
<< viali >>
rect -746 1027 2144 1086
rect -746 994 -715 1027
rect -715 994 2144 1027
<< metal1 >>
rect -888 1160 2204 1176
rect -888 1086 2208 1160
rect -888 994 -746 1086
rect 2144 994 2208 1086
rect -888 958 2208 994
rect -616 -202 -570 -12
rect 700 -214 746 -22
rect 2016 -200 2062 -44
use sky130_fd_pr__pfet_g5v0d10v5_8ZATBS  sky130_fd_pr__pfet_g5v0d10v5_8ZATBS_0
timestamp 1738973041
transform -1 0 -264 0 1 214
box -424 -336 424 252
use sky130_fd_pr__pfet_g5v0d10v5_8ZATBS  sky130_fd_pr__pfet_g5v0d10v5_8ZATBS_1
timestamp 1738973041
transform 1 0 1710 0 1 214
box -424 -336 424 252
use sky130_fd_pr__pfet_g5v0d10v5_8ZATBS  sky130_fd_pr__pfet_g5v0d10v5_8ZATBS_2
timestamp 1738973041
transform -1 0 -264 0 1 682
box -424 -336 424 252
use sky130_fd_pr__pfet_g5v0d10v5_8ZATBS  sky130_fd_pr__pfet_g5v0d10v5_8ZATBS_3
timestamp 1738973041
transform 1 0 1710 0 1 682
box -424 -336 424 252
use sky130_fd_pr__pfet_g5v0d10v5_ALBTBJ  sky130_fd_pr__pfet_g5v0d10v5_ALBTBJ_1
timestamp 1738973041
transform 1 0 723 0 1 214
box -753 -282 859 372
use sky130_fd_pr__pfet_g5v0d10v5_ALBTBJ  sky130_fd_pr__pfet_g5v0d10v5_ALBTBJ_2
timestamp 1738973041
transform 1 0 723 0 1 682
box -753 -282 859 372
<< labels >>
flabel metal1 -868 1022 -814 1136 0 FreeSans 1600 0 0 0 VDD
port 1 nsew
flabel metal1 710 -194 740 -168 0 FreeSans 1600 0 0 0 IB
port 4 nsew
flabel metal1 -610 -190 -580 -166 0 FreeSans 1600 0 0 0 IA
port 6 nsew
<< end >>
