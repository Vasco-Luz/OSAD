magic
tech sky130A
magscale 1 2
timestamp 1743851084
<< pwell >>
rect -26 -26 108 1106
<< psubdiff >>
rect 0 1033 82 1080
rect 0 999 24 1033
rect 58 999 82 1033
rect 0 965 82 999
rect 0 931 24 965
rect 58 931 82 965
rect 0 897 82 931
rect 0 863 24 897
rect 58 863 82 897
rect 0 829 82 863
rect 0 795 24 829
rect 58 795 82 829
rect 0 761 82 795
rect 0 727 24 761
rect 58 727 82 761
rect 0 693 82 727
rect 0 659 24 693
rect 58 659 82 693
rect 0 625 82 659
rect 0 591 24 625
rect 58 591 82 625
rect 0 557 82 591
rect 0 523 24 557
rect 58 523 82 557
rect 0 489 82 523
rect 0 455 24 489
rect 58 455 82 489
rect 0 421 82 455
rect 0 387 24 421
rect 58 387 82 421
rect 0 353 82 387
rect 0 319 24 353
rect 58 319 82 353
rect 0 285 82 319
rect 0 251 24 285
rect 58 251 82 285
rect 0 217 82 251
rect 0 183 24 217
rect 58 183 82 217
rect 0 149 82 183
rect 0 115 24 149
rect 58 115 82 149
rect 0 81 82 115
rect 0 47 24 81
rect 58 47 82 81
rect 0 0 82 47
<< psubdiffcont >>
rect 24 999 58 1033
rect 24 931 58 965
rect 24 863 58 897
rect 24 795 58 829
rect 24 727 58 761
rect 24 659 58 693
rect 24 591 58 625
rect 24 523 58 557
rect 24 455 58 489
rect 24 387 58 421
rect 24 319 58 353
rect 24 251 58 285
rect 24 183 58 217
rect 24 115 58 149
rect 24 47 58 81
<< locali >>
rect 0 1033 82 1080
rect 0 999 24 1033
rect 58 999 82 1033
rect 0 965 82 999
rect 0 931 24 965
rect 58 931 82 965
rect 0 897 82 931
rect 0 863 24 897
rect 58 863 82 897
rect 0 829 82 863
rect 0 795 24 829
rect 58 795 82 829
rect 0 761 82 795
rect 0 727 24 761
rect 58 727 82 761
rect 0 693 82 727
rect 0 659 24 693
rect 58 659 82 693
rect 0 625 82 659
rect 0 591 24 625
rect 58 591 82 625
rect 0 557 82 591
rect 0 523 24 557
rect 58 523 82 557
rect 0 489 82 523
rect 0 455 24 489
rect 58 455 82 489
rect 0 421 82 455
rect 0 387 24 421
rect 58 387 82 421
rect 0 353 82 387
rect 0 319 24 353
rect 58 319 82 353
rect 0 285 82 319
rect 0 251 24 285
rect 58 251 82 285
rect 0 217 82 251
rect 0 183 24 217
rect 58 183 82 217
rect 0 149 82 183
rect 0 115 24 149
rect 58 115 82 149
rect 0 81 82 115
rect 0 47 24 81
rect 58 47 82 81
rect 0 0 82 47
<< end >>
