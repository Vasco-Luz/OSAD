** sch_path:
*+ /home/vasco/Desktop/sky130A/amplifiers/single_stage_amps/basic_stages/cs_resistor_stage/genetic_automatic/cs_resistor_stage_test.sch
**.subckt cs_resistor_stage_test
Vmeas VDD net1 0
.save i(vmeas)
V1 VDD GND VDD
.save i(v1)
V2 net2 GND vin
.save i(v2)
R2 VOUT GND 10G m=1
XR6 VOUT net1 VDD sky130_fd_pr__res_high_po_0p35 L=R1 mult=2 m=2
V4 VIN net2 ac 1.0 sin (0 100u 100k)
.save i(v4)
XM5 VOUT VIN GND GND sky130_fd_pr__nfet_g5v0d10v5 L=L1 W=W1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
**** begin user architecture code

**************************************************************
**************************************************************
**************************************************************
**************************************************************
**************************************************************
*LIBs*********************************************************
**************************************************************
**************************************************************
**************************************************************
**************************************************************
**************************************************************
*.lib /home/vasco/Desktop/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
* chose the corners in the corner file
* tt_mm for mismatch
* ss ff sf fs standart corners
* ll hh lh hl capacitor and resistors corners
* mc for total process variation including corners
**************************************************************
**************************************************************
**************************************************************
**************************************************************
**************************************************************
*Corners/montecarlo options***********************************
**************************************************************
**************************************************************
**************************************************************
**************************************************************
**************************************************************
.TEMP 27
**************************************************************
**************************************************************
**************************************************************
**************************************************************
*SIMULATION and Plots*****************************************
**************************************************************
**************************************************************
**************************************************************
**************************************************************


.control
.param R1 = 5
.param L1 = 0.5
.param VDD = 5
.param W1 = 50
.param vin =  2



save all




.endc


.param mc_mm_switch=0
.param mc_pr_switch=0
.include /home/vasco/Desktop/pdk/sky130A/libs.tech/ngspice/corners/tt.spice
.include /home/vasco/Desktop/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/vasco/Desktop/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/vasco/Desktop/pdk/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends
.GLOBAL GND
.end
