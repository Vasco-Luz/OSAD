magic
tech sky130A
magscale 1 2
timestamp 1740488682
<< metal3 >>
rect -2092 1772 -120 1800
rect -2092 148 -204 1772
rect -140 148 -120 1772
rect -2092 120 -120 148
rect 120 1772 2092 1800
rect 120 148 2008 1772
rect 2072 148 2092 1772
rect 120 120 2092 148
rect -2092 -148 -120 -120
rect -2092 -1772 -204 -148
rect -140 -1772 -120 -148
rect -2092 -1800 -120 -1772
rect 120 -148 2092 -120
rect 120 -1772 2008 -148
rect 2072 -1772 2092 -148
rect 120 -1800 2092 -1772
<< via3 >>
rect -204 148 -140 1772
rect 2008 148 2072 1772
rect -204 -1772 -140 -148
rect 2008 -1772 2072 -148
<< mimcap >>
rect -2052 1720 -452 1760
rect -2052 200 -2012 1720
rect -492 200 -452 1720
rect -2052 160 -452 200
rect 160 1720 1760 1760
rect 160 200 200 1720
rect 1720 200 1760 1720
rect 160 160 1760 200
rect -2052 -200 -452 -160
rect -2052 -1720 -2012 -200
rect -492 -1720 -452 -200
rect -2052 -1760 -452 -1720
rect 160 -200 1760 -160
rect 160 -1720 200 -200
rect 1720 -1720 1760 -200
rect 160 -1760 1760 -1720
<< mimcapcontact >>
rect -2012 200 -492 1720
rect 200 200 1720 1720
rect -2012 -1720 -492 -200
rect 200 -1720 1720 -200
<< metal4 >>
rect -1304 1721 -1200 1920
rect -224 1772 -120 1920
rect -2013 1720 -491 1721
rect -2013 200 -2012 1720
rect -492 200 -491 1720
rect -2013 199 -491 200
rect -1304 -199 -1200 199
rect -224 148 -204 1772
rect -140 148 -120 1772
rect 908 1721 1012 1920
rect 1988 1772 2092 1920
rect 199 1720 1721 1721
rect 199 200 200 1720
rect 1720 200 1721 1720
rect 199 199 1721 200
rect -224 -148 -120 148
rect -2013 -200 -491 -199
rect -2013 -1720 -2012 -200
rect -492 -1720 -491 -200
rect -2013 -1721 -491 -1720
rect -1304 -1920 -1200 -1721
rect -224 -1772 -204 -148
rect -140 -1772 -120 -148
rect 908 -199 1012 199
rect 1988 148 2008 1772
rect 2072 148 2092 1772
rect 1988 -148 2092 148
rect 199 -200 1721 -199
rect 199 -1720 200 -200
rect 1720 -1720 1721 -200
rect 199 -1721 1721 -1720
rect -224 -1920 -120 -1772
rect 908 -1920 1012 -1721
rect 1988 -1772 2008 -148
rect 2072 -1772 2092 -148
rect 1988 -1920 2092 -1772
<< properties >>
string FIXED_BBOX 120 120 1800 1800
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 8 l 8 val 134.08 carea 2.00 cperi 0.19 class capacitor nx 2 ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
