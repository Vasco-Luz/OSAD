magic
tech sky130A
magscale 1 2
timestamp 1740488222
<< metal3 >>
rect -892 572 -120 600
rect -892 148 -204 572
rect -140 148 -120 572
rect -892 120 -120 148
rect 120 572 892 600
rect 120 148 808 572
rect 872 148 892 572
rect 120 120 892 148
rect -892 -148 -120 -120
rect -892 -572 -204 -148
rect -140 -572 -120 -148
rect -892 -600 -120 -572
rect 120 -148 892 -120
rect 120 -572 808 -148
rect 872 -572 892 -148
rect 120 -600 892 -572
<< via3 >>
rect -204 148 -140 572
rect 808 148 872 572
rect -204 -572 -140 -148
rect 808 -572 872 -148
<< mimcap >>
rect -852 520 -452 560
rect -852 200 -812 520
rect -492 200 -452 520
rect -852 160 -452 200
rect 160 520 560 560
rect 160 200 200 520
rect 520 200 560 520
rect 160 160 560 200
rect -852 -200 -452 -160
rect -852 -520 -812 -200
rect -492 -520 -452 -200
rect -852 -560 -452 -520
rect 160 -200 560 -160
rect 160 -520 200 -200
rect 520 -520 560 -200
rect 160 -560 560 -520
<< mimcapcontact >>
rect -812 200 -492 520
rect 200 200 520 520
rect -812 -520 -492 -200
rect 200 -520 520 -200
<< metal4 >>
rect -704 521 -600 720
rect -224 572 -120 720
rect -813 520 -491 521
rect -813 200 -812 520
rect -492 200 -491 520
rect -813 199 -491 200
rect -704 -199 -600 199
rect -224 148 -204 572
rect -140 148 -120 572
rect 308 521 412 720
rect 788 572 892 720
rect 199 520 521 521
rect 199 200 200 520
rect 520 200 521 520
rect 199 199 521 200
rect -224 -148 -120 148
rect -813 -200 -491 -199
rect -813 -520 -812 -200
rect -492 -520 -491 -200
rect -813 -521 -491 -520
rect -704 -720 -600 -521
rect -224 -572 -204 -148
rect -140 -572 -120 -148
rect 308 -199 412 199
rect 788 148 808 572
rect 872 148 892 572
rect 788 -148 892 148
rect 199 -200 521 -199
rect 199 -520 200 -200
rect 520 -520 521 -200
rect 199 -521 521 -520
rect -224 -720 -120 -572
rect 308 -720 412 -521
rect 788 -572 808 -148
rect 872 -572 892 -148
rect 788 -720 892 -572
<< properties >>
string FIXED_BBOX 120 120 600 600
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.0 l 2.0 val 9.52 carea 2.00 cperi 0.19 class capacitor nx 2 ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
