** sch_path: /foss/designs/OSAD/my_ip/LIB/ihp-sg13g2/FD_opamp001/first_stage.sch
**.subckt first_stage VDD VSS VB VIN+ VIN- VOUT- VOUT+ VB2 VCM V_COMP+ V_COMP-
*.iopin VDD
*.iopin VSS
*.iopin VB
*.iopin VIN+
*.iopin VIN-
*.iopin VOUT-
*.iopin VOUT+
*.iopin VB2
*.iopin VCM
*.iopin V_COMP+
*.iopin V_COMP-
XM13 net2 VB VSS VSS sg13_hv_nmos w=4.5u l=2u ng=2 m=2
XM14 net1 VCM net3 VSS sg13_hv_nmos w=5u l=1.5u ng=2 m=2
XM15 VB2 VCM net1 VSS sg13_hv_nmos w=5u l=1.5u ng=2 m=2
XM16 VB2 VB2 VDD VDD sg13_hv_pmos w=2.2u l=3u ng=2 m=2
Vmeas2 net3 net2 0
.save i(vmeas2)
XM17 V_COMP+ VIN+ net4 VSS sg13_hv_nmos w=5u l=1.5u ng=2 m=2
XM18 VOUT- VIN+ V_COMP+ VSS sg13_hv_nmos w=5u l=1.5u ng=2 m=2
XM19 V_COMP- VIN- net4 VSS sg13_hv_nmos w=5u l=1.5u ng=2 m=2
XM20 VOUT+ VIN- V_COMP- VSS sg13_hv_nmos w=5u l=1.5u ng=2 m=2
XM21 net4 VB VSS VSS sg13_hv_nmos w=4.5u l=2u ng=2 m=2
XM22 net4 VB VSS VSS sg13_hv_nmos w=4.5u l=2u ng=2 m=2
XM23 VOUT+ VB2 VDD VDD sg13_hv_pmos w=2.2u l=3u ng=2 m=2
XM24 VOUT- VB2 VDD VDD sg13_hv_pmos w=2.2u l=3u ng=2 m=2
**.ends
.end
