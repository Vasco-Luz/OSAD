magic
tech sky130A
magscale 1 2
timestamp 1693698878
<< nwell >>
rect -883 -1297 883 1297
<< mvpmos >>
rect -625 -1000 -465 1000
rect -407 -1000 -247 1000
rect -189 -1000 -29 1000
rect 29 -1000 189 1000
rect 247 -1000 407 1000
rect 465 -1000 625 1000
<< mvpdiff >>
rect -683 988 -625 1000
rect -683 -988 -671 988
rect -637 -988 -625 988
rect -683 -1000 -625 -988
rect -465 988 -407 1000
rect -465 -988 -453 988
rect -419 -988 -407 988
rect -465 -1000 -407 -988
rect -247 988 -189 1000
rect -247 -988 -235 988
rect -201 -988 -189 988
rect -247 -1000 -189 -988
rect -29 988 29 1000
rect -29 -988 -17 988
rect 17 -988 29 988
rect -29 -1000 29 -988
rect 189 988 247 1000
rect 189 -988 201 988
rect 235 -988 247 988
rect 189 -1000 247 -988
rect 407 988 465 1000
rect 407 -988 419 988
rect 453 -988 465 988
rect 407 -1000 465 -988
rect 625 988 683 1000
rect 625 -988 637 988
rect 671 -988 683 988
rect 625 -1000 683 -988
<< mvpdiffc >>
rect -671 -988 -637 988
rect -453 -988 -419 988
rect -235 -988 -201 988
rect -17 -988 17 988
rect 201 -988 235 988
rect 419 -988 453 988
rect 637 -988 671 988
<< mvnsubdiff >>
rect -817 1219 817 1231
rect -817 1185 -709 1219
rect 709 1185 817 1219
rect -817 1173 817 1185
rect -817 1123 -759 1173
rect -817 -1123 -805 1123
rect -771 -1123 -759 1123
rect 759 1123 817 1173
rect -817 -1173 -759 -1123
rect 759 -1123 771 1123
rect 805 -1123 817 1123
rect 759 -1173 817 -1123
rect -817 -1185 817 -1173
rect -817 -1219 -709 -1185
rect 709 -1219 817 -1185
rect -817 -1231 817 -1219
<< mvnsubdiffcont >>
rect -709 1185 709 1219
rect -805 -1123 -771 1123
rect 771 -1123 805 1123
rect -709 -1219 709 -1185
<< poly >>
rect -625 1081 -465 1097
rect -625 1047 -609 1081
rect -481 1047 -465 1081
rect -625 1000 -465 1047
rect -407 1081 -247 1097
rect -407 1047 -391 1081
rect -263 1047 -247 1081
rect -407 1000 -247 1047
rect -189 1081 -29 1097
rect -189 1047 -173 1081
rect -45 1047 -29 1081
rect -189 1000 -29 1047
rect 29 1081 189 1097
rect 29 1047 45 1081
rect 173 1047 189 1081
rect 29 1000 189 1047
rect 247 1081 407 1097
rect 247 1047 263 1081
rect 391 1047 407 1081
rect 247 1000 407 1047
rect 465 1081 625 1097
rect 465 1047 481 1081
rect 609 1047 625 1081
rect 465 1000 625 1047
rect -625 -1047 -465 -1000
rect -625 -1081 -609 -1047
rect -481 -1081 -465 -1047
rect -625 -1097 -465 -1081
rect -407 -1047 -247 -1000
rect -407 -1081 -391 -1047
rect -263 -1081 -247 -1047
rect -407 -1097 -247 -1081
rect -189 -1047 -29 -1000
rect -189 -1081 -173 -1047
rect -45 -1081 -29 -1047
rect -189 -1097 -29 -1081
rect 29 -1047 189 -1000
rect 29 -1081 45 -1047
rect 173 -1081 189 -1047
rect 29 -1097 189 -1081
rect 247 -1047 407 -1000
rect 247 -1081 263 -1047
rect 391 -1081 407 -1047
rect 247 -1097 407 -1081
rect 465 -1047 625 -1000
rect 465 -1081 481 -1047
rect 609 -1081 625 -1047
rect 465 -1097 625 -1081
<< polycont >>
rect -609 1047 -481 1081
rect -391 1047 -263 1081
rect -173 1047 -45 1081
rect 45 1047 173 1081
rect 263 1047 391 1081
rect 481 1047 609 1081
rect -609 -1081 -481 -1047
rect -391 -1081 -263 -1047
rect -173 -1081 -45 -1047
rect 45 -1081 173 -1047
rect 263 -1081 391 -1047
rect 481 -1081 609 -1047
<< locali >>
rect -805 1185 -709 1219
rect 709 1185 805 1219
rect -805 1123 -771 1185
rect 771 1123 805 1185
rect -625 1047 -609 1081
rect -481 1047 -465 1081
rect -407 1047 -391 1081
rect -263 1047 -247 1081
rect -189 1047 -173 1081
rect -45 1047 -29 1081
rect 29 1047 45 1081
rect 173 1047 189 1081
rect 247 1047 263 1081
rect 391 1047 407 1081
rect 465 1047 481 1081
rect 609 1047 625 1081
rect -671 988 -637 1004
rect -671 -1004 -637 -988
rect -453 988 -419 1004
rect -453 -1004 -419 -988
rect -235 988 -201 1004
rect -235 -1004 -201 -988
rect -17 988 17 1004
rect -17 -1004 17 -988
rect 201 988 235 1004
rect 201 -1004 235 -988
rect 419 988 453 1004
rect 419 -1004 453 -988
rect 637 988 671 1004
rect 637 -1004 671 -988
rect -625 -1081 -609 -1047
rect -481 -1081 -465 -1047
rect -407 -1081 -391 -1047
rect -263 -1081 -247 -1047
rect -189 -1081 -173 -1047
rect -45 -1081 -29 -1047
rect 29 -1081 45 -1047
rect 173 -1081 189 -1047
rect 247 -1081 263 -1047
rect 391 -1081 407 -1047
rect 465 -1081 481 -1047
rect 609 -1081 625 -1047
rect -805 -1185 -771 -1123
rect 771 -1185 805 -1123
rect -805 -1219 -709 -1185
rect 709 -1219 805 -1185
<< viali >>
rect -609 1047 -481 1081
rect -391 1047 -263 1081
rect -173 1047 -45 1081
rect 45 1047 173 1081
rect 263 1047 391 1081
rect 481 1047 609 1081
rect -671 -988 -637 988
rect -453 -988 -419 988
rect -235 -988 -201 988
rect -17 -988 17 988
rect 201 -988 235 988
rect 419 -988 453 988
rect 637 -988 671 988
rect -609 -1081 -481 -1047
rect -391 -1081 -263 -1047
rect -173 -1081 -45 -1047
rect 45 -1081 173 -1047
rect 263 -1081 391 -1047
rect 481 -1081 609 -1047
<< metal1 >>
rect -621 1081 -469 1087
rect -621 1047 -609 1081
rect -481 1047 -469 1081
rect -621 1041 -469 1047
rect -403 1081 -251 1087
rect -403 1047 -391 1081
rect -263 1047 -251 1081
rect -403 1041 -251 1047
rect -185 1081 -33 1087
rect -185 1047 -173 1081
rect -45 1047 -33 1081
rect -185 1041 -33 1047
rect 33 1081 185 1087
rect 33 1047 45 1081
rect 173 1047 185 1081
rect 33 1041 185 1047
rect 251 1081 403 1087
rect 251 1047 263 1081
rect 391 1047 403 1081
rect 251 1041 403 1047
rect 469 1081 621 1087
rect 469 1047 481 1081
rect 609 1047 621 1081
rect 469 1041 621 1047
rect -677 988 -631 1000
rect -677 -988 -671 988
rect -637 -988 -631 988
rect -677 -1000 -631 -988
rect -459 988 -413 1000
rect -459 -988 -453 988
rect -419 -988 -413 988
rect -459 -1000 -413 -988
rect -241 988 -195 1000
rect -241 -988 -235 988
rect -201 -988 -195 988
rect -241 -1000 -195 -988
rect -23 988 23 1000
rect -23 -988 -17 988
rect 17 -988 23 988
rect -23 -1000 23 -988
rect 195 988 241 1000
rect 195 -988 201 988
rect 235 -988 241 988
rect 195 -1000 241 -988
rect 413 988 459 1000
rect 413 -988 419 988
rect 453 -988 459 988
rect 413 -1000 459 -988
rect 631 988 677 1000
rect 631 -988 637 988
rect 671 -988 677 988
rect 631 -1000 677 -988
rect -621 -1047 -469 -1041
rect -621 -1081 -609 -1047
rect -481 -1081 -469 -1047
rect -621 -1087 -469 -1081
rect -403 -1047 -251 -1041
rect -403 -1081 -391 -1047
rect -263 -1081 -251 -1047
rect -403 -1087 -251 -1081
rect -185 -1047 -33 -1041
rect -185 -1081 -173 -1047
rect -45 -1081 -33 -1047
rect -185 -1087 -33 -1081
rect 33 -1047 185 -1041
rect 33 -1081 45 -1047
rect 173 -1081 185 -1047
rect 33 -1087 185 -1081
rect 251 -1047 403 -1041
rect 251 -1081 263 -1047
rect 391 -1081 403 -1047
rect 251 -1087 403 -1081
rect 469 -1047 621 -1041
rect 469 -1081 481 -1047
rect 609 -1081 621 -1047
rect 469 -1087 621 -1081
<< properties >>
string FIXED_BBOX -788 -1202 788 1202
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 10 l 0.8 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
