magic
tech sky130A
magscale 1 2
timestamp 1743851084
<< pwell >>
rect -26 -26 108 13026
<< psubdiff >>
rect 0 12977 82 13000
rect 0 12943 24 12977
rect 58 12943 82 12977
rect 0 12909 82 12943
rect 0 12875 24 12909
rect 58 12875 82 12909
rect 0 12841 82 12875
rect 0 12807 24 12841
rect 58 12807 82 12841
rect 0 12773 82 12807
rect 0 12739 24 12773
rect 58 12739 82 12773
rect 0 12705 82 12739
rect 0 12671 24 12705
rect 58 12671 82 12705
rect 0 12637 82 12671
rect 0 12603 24 12637
rect 58 12603 82 12637
rect 0 12569 82 12603
rect 0 12535 24 12569
rect 58 12535 82 12569
rect 0 12501 82 12535
rect 0 12467 24 12501
rect 58 12467 82 12501
rect 0 12433 82 12467
rect 0 12399 24 12433
rect 58 12399 82 12433
rect 0 12365 82 12399
rect 0 12331 24 12365
rect 58 12331 82 12365
rect 0 12297 82 12331
rect 0 12263 24 12297
rect 58 12263 82 12297
rect 0 12229 82 12263
rect 0 12195 24 12229
rect 58 12195 82 12229
rect 0 12161 82 12195
rect 0 12127 24 12161
rect 58 12127 82 12161
rect 0 12093 82 12127
rect 0 12059 24 12093
rect 58 12059 82 12093
rect 0 12025 82 12059
rect 0 11991 24 12025
rect 58 11991 82 12025
rect 0 11957 82 11991
rect 0 11923 24 11957
rect 58 11923 82 11957
rect 0 11889 82 11923
rect 0 11855 24 11889
rect 58 11855 82 11889
rect 0 11821 82 11855
rect 0 11787 24 11821
rect 58 11787 82 11821
rect 0 11753 82 11787
rect 0 11719 24 11753
rect 58 11719 82 11753
rect 0 11685 82 11719
rect 0 11651 24 11685
rect 58 11651 82 11685
rect 0 11617 82 11651
rect 0 11583 24 11617
rect 58 11583 82 11617
rect 0 11549 82 11583
rect 0 11515 24 11549
rect 58 11515 82 11549
rect 0 11481 82 11515
rect 0 11447 24 11481
rect 58 11447 82 11481
rect 0 11413 82 11447
rect 0 11379 24 11413
rect 58 11379 82 11413
rect 0 11345 82 11379
rect 0 11311 24 11345
rect 58 11311 82 11345
rect 0 11277 82 11311
rect 0 11243 24 11277
rect 58 11243 82 11277
rect 0 11209 82 11243
rect 0 11175 24 11209
rect 58 11175 82 11209
rect 0 11141 82 11175
rect 0 11107 24 11141
rect 58 11107 82 11141
rect 0 11073 82 11107
rect 0 11039 24 11073
rect 58 11039 82 11073
rect 0 11005 82 11039
rect 0 10971 24 11005
rect 58 10971 82 11005
rect 0 10937 82 10971
rect 0 10903 24 10937
rect 58 10903 82 10937
rect 0 10869 82 10903
rect 0 10835 24 10869
rect 58 10835 82 10869
rect 0 10801 82 10835
rect 0 10767 24 10801
rect 58 10767 82 10801
rect 0 10733 82 10767
rect 0 10699 24 10733
rect 58 10699 82 10733
rect 0 10665 82 10699
rect 0 10631 24 10665
rect 58 10631 82 10665
rect 0 10597 82 10631
rect 0 10563 24 10597
rect 58 10563 82 10597
rect 0 10529 82 10563
rect 0 10495 24 10529
rect 58 10495 82 10529
rect 0 10461 82 10495
rect 0 10427 24 10461
rect 58 10427 82 10461
rect 0 10393 82 10427
rect 0 10359 24 10393
rect 58 10359 82 10393
rect 0 10325 82 10359
rect 0 10291 24 10325
rect 58 10291 82 10325
rect 0 10257 82 10291
rect 0 10223 24 10257
rect 58 10223 82 10257
rect 0 10189 82 10223
rect 0 10155 24 10189
rect 58 10155 82 10189
rect 0 10121 82 10155
rect 0 10087 24 10121
rect 58 10087 82 10121
rect 0 10053 82 10087
rect 0 10019 24 10053
rect 58 10019 82 10053
rect 0 9985 82 10019
rect 0 9951 24 9985
rect 58 9951 82 9985
rect 0 9917 82 9951
rect 0 9883 24 9917
rect 58 9883 82 9917
rect 0 9849 82 9883
rect 0 9815 24 9849
rect 58 9815 82 9849
rect 0 9781 82 9815
rect 0 9747 24 9781
rect 58 9747 82 9781
rect 0 9713 82 9747
rect 0 9679 24 9713
rect 58 9679 82 9713
rect 0 9645 82 9679
rect 0 9611 24 9645
rect 58 9611 82 9645
rect 0 9577 82 9611
rect 0 9543 24 9577
rect 58 9543 82 9577
rect 0 9509 82 9543
rect 0 9475 24 9509
rect 58 9475 82 9509
rect 0 9441 82 9475
rect 0 9407 24 9441
rect 58 9407 82 9441
rect 0 9373 82 9407
rect 0 9339 24 9373
rect 58 9339 82 9373
rect 0 9305 82 9339
rect 0 9271 24 9305
rect 58 9271 82 9305
rect 0 9237 82 9271
rect 0 9203 24 9237
rect 58 9203 82 9237
rect 0 9169 82 9203
rect 0 9135 24 9169
rect 58 9135 82 9169
rect 0 9101 82 9135
rect 0 9067 24 9101
rect 58 9067 82 9101
rect 0 9033 82 9067
rect 0 8999 24 9033
rect 58 8999 82 9033
rect 0 8965 82 8999
rect 0 8931 24 8965
rect 58 8931 82 8965
rect 0 8897 82 8931
rect 0 8863 24 8897
rect 58 8863 82 8897
rect 0 8829 82 8863
rect 0 8795 24 8829
rect 58 8795 82 8829
rect 0 8761 82 8795
rect 0 8727 24 8761
rect 58 8727 82 8761
rect 0 8693 82 8727
rect 0 8659 24 8693
rect 58 8659 82 8693
rect 0 8625 82 8659
rect 0 8591 24 8625
rect 58 8591 82 8625
rect 0 8557 82 8591
rect 0 8523 24 8557
rect 58 8523 82 8557
rect 0 8489 82 8523
rect 0 8455 24 8489
rect 58 8455 82 8489
rect 0 8421 82 8455
rect 0 8387 24 8421
rect 58 8387 82 8421
rect 0 8353 82 8387
rect 0 8319 24 8353
rect 58 8319 82 8353
rect 0 8285 82 8319
rect 0 8251 24 8285
rect 58 8251 82 8285
rect 0 8217 82 8251
rect 0 8183 24 8217
rect 58 8183 82 8217
rect 0 8149 82 8183
rect 0 8115 24 8149
rect 58 8115 82 8149
rect 0 8081 82 8115
rect 0 8047 24 8081
rect 58 8047 82 8081
rect 0 8013 82 8047
rect 0 7979 24 8013
rect 58 7979 82 8013
rect 0 7945 82 7979
rect 0 7911 24 7945
rect 58 7911 82 7945
rect 0 7877 82 7911
rect 0 7843 24 7877
rect 58 7843 82 7877
rect 0 7809 82 7843
rect 0 7775 24 7809
rect 58 7775 82 7809
rect 0 7741 82 7775
rect 0 7707 24 7741
rect 58 7707 82 7741
rect 0 7673 82 7707
rect 0 7639 24 7673
rect 58 7639 82 7673
rect 0 7605 82 7639
rect 0 7571 24 7605
rect 58 7571 82 7605
rect 0 7537 82 7571
rect 0 7503 24 7537
rect 58 7503 82 7537
rect 0 7469 82 7503
rect 0 7435 24 7469
rect 58 7435 82 7469
rect 0 7401 82 7435
rect 0 7367 24 7401
rect 58 7367 82 7401
rect 0 7333 82 7367
rect 0 7299 24 7333
rect 58 7299 82 7333
rect 0 7265 82 7299
rect 0 7231 24 7265
rect 58 7231 82 7265
rect 0 7197 82 7231
rect 0 7163 24 7197
rect 58 7163 82 7197
rect 0 7129 82 7163
rect 0 7095 24 7129
rect 58 7095 82 7129
rect 0 7061 82 7095
rect 0 7027 24 7061
rect 58 7027 82 7061
rect 0 6993 82 7027
rect 0 6959 24 6993
rect 58 6959 82 6993
rect 0 6925 82 6959
rect 0 6891 24 6925
rect 58 6891 82 6925
rect 0 6857 82 6891
rect 0 6823 24 6857
rect 58 6823 82 6857
rect 0 6789 82 6823
rect 0 6755 24 6789
rect 58 6755 82 6789
rect 0 6721 82 6755
rect 0 6687 24 6721
rect 58 6687 82 6721
rect 0 6653 82 6687
rect 0 6619 24 6653
rect 58 6619 82 6653
rect 0 6585 82 6619
rect 0 6551 24 6585
rect 58 6551 82 6585
rect 0 6517 82 6551
rect 0 6483 24 6517
rect 58 6483 82 6517
rect 0 6449 82 6483
rect 0 6415 24 6449
rect 58 6415 82 6449
rect 0 6381 82 6415
rect 0 6347 24 6381
rect 58 6347 82 6381
rect 0 6313 82 6347
rect 0 6279 24 6313
rect 58 6279 82 6313
rect 0 6245 82 6279
rect 0 6211 24 6245
rect 58 6211 82 6245
rect 0 6177 82 6211
rect 0 6143 24 6177
rect 58 6143 82 6177
rect 0 6109 82 6143
rect 0 6075 24 6109
rect 58 6075 82 6109
rect 0 6041 82 6075
rect 0 6007 24 6041
rect 58 6007 82 6041
rect 0 5973 82 6007
rect 0 5939 24 5973
rect 58 5939 82 5973
rect 0 5905 82 5939
rect 0 5871 24 5905
rect 58 5871 82 5905
rect 0 5837 82 5871
rect 0 5803 24 5837
rect 58 5803 82 5837
rect 0 5769 82 5803
rect 0 5735 24 5769
rect 58 5735 82 5769
rect 0 5701 82 5735
rect 0 5667 24 5701
rect 58 5667 82 5701
rect 0 5633 82 5667
rect 0 5599 24 5633
rect 58 5599 82 5633
rect 0 5565 82 5599
rect 0 5531 24 5565
rect 58 5531 82 5565
rect 0 5497 82 5531
rect 0 5463 24 5497
rect 58 5463 82 5497
rect 0 5429 82 5463
rect 0 5395 24 5429
rect 58 5395 82 5429
rect 0 5361 82 5395
rect 0 5327 24 5361
rect 58 5327 82 5361
rect 0 5293 82 5327
rect 0 5259 24 5293
rect 58 5259 82 5293
rect 0 5225 82 5259
rect 0 5191 24 5225
rect 58 5191 82 5225
rect 0 5157 82 5191
rect 0 5123 24 5157
rect 58 5123 82 5157
rect 0 5089 82 5123
rect 0 5055 24 5089
rect 58 5055 82 5089
rect 0 5021 82 5055
rect 0 4987 24 5021
rect 58 4987 82 5021
rect 0 4953 82 4987
rect 0 4919 24 4953
rect 58 4919 82 4953
rect 0 4885 82 4919
rect 0 4851 24 4885
rect 58 4851 82 4885
rect 0 4817 82 4851
rect 0 4783 24 4817
rect 58 4783 82 4817
rect 0 4749 82 4783
rect 0 4715 24 4749
rect 58 4715 82 4749
rect 0 4681 82 4715
rect 0 4647 24 4681
rect 58 4647 82 4681
rect 0 4613 82 4647
rect 0 4579 24 4613
rect 58 4579 82 4613
rect 0 4545 82 4579
rect 0 4511 24 4545
rect 58 4511 82 4545
rect 0 4477 82 4511
rect 0 4443 24 4477
rect 58 4443 82 4477
rect 0 4409 82 4443
rect 0 4375 24 4409
rect 58 4375 82 4409
rect 0 4341 82 4375
rect 0 4307 24 4341
rect 58 4307 82 4341
rect 0 4273 82 4307
rect 0 4239 24 4273
rect 58 4239 82 4273
rect 0 4205 82 4239
rect 0 4171 24 4205
rect 58 4171 82 4205
rect 0 4137 82 4171
rect 0 4103 24 4137
rect 58 4103 82 4137
rect 0 4069 82 4103
rect 0 4035 24 4069
rect 58 4035 82 4069
rect 0 4001 82 4035
rect 0 3967 24 4001
rect 58 3967 82 4001
rect 0 3933 82 3967
rect 0 3899 24 3933
rect 58 3899 82 3933
rect 0 3865 82 3899
rect 0 3831 24 3865
rect 58 3831 82 3865
rect 0 3797 82 3831
rect 0 3763 24 3797
rect 58 3763 82 3797
rect 0 3729 82 3763
rect 0 3695 24 3729
rect 58 3695 82 3729
rect 0 3661 82 3695
rect 0 3627 24 3661
rect 58 3627 82 3661
rect 0 3593 82 3627
rect 0 3559 24 3593
rect 58 3559 82 3593
rect 0 3525 82 3559
rect 0 3491 24 3525
rect 58 3491 82 3525
rect 0 3457 82 3491
rect 0 3423 24 3457
rect 58 3423 82 3457
rect 0 3389 82 3423
rect 0 3355 24 3389
rect 58 3355 82 3389
rect 0 3321 82 3355
rect 0 3287 24 3321
rect 58 3287 82 3321
rect 0 3253 82 3287
rect 0 3219 24 3253
rect 58 3219 82 3253
rect 0 3185 82 3219
rect 0 3151 24 3185
rect 58 3151 82 3185
rect 0 3117 82 3151
rect 0 3083 24 3117
rect 58 3083 82 3117
rect 0 3049 82 3083
rect 0 3015 24 3049
rect 58 3015 82 3049
rect 0 2981 82 3015
rect 0 2947 24 2981
rect 58 2947 82 2981
rect 0 2913 82 2947
rect 0 2879 24 2913
rect 58 2879 82 2913
rect 0 2845 82 2879
rect 0 2811 24 2845
rect 58 2811 82 2845
rect 0 2777 82 2811
rect 0 2743 24 2777
rect 58 2743 82 2777
rect 0 2709 82 2743
rect 0 2675 24 2709
rect 58 2675 82 2709
rect 0 2641 82 2675
rect 0 2607 24 2641
rect 58 2607 82 2641
rect 0 2573 82 2607
rect 0 2539 24 2573
rect 58 2539 82 2573
rect 0 2505 82 2539
rect 0 2471 24 2505
rect 58 2471 82 2505
rect 0 2437 82 2471
rect 0 2403 24 2437
rect 58 2403 82 2437
rect 0 2369 82 2403
rect 0 2335 24 2369
rect 58 2335 82 2369
rect 0 2301 82 2335
rect 0 2267 24 2301
rect 58 2267 82 2301
rect 0 2233 82 2267
rect 0 2199 24 2233
rect 58 2199 82 2233
rect 0 2165 82 2199
rect 0 2131 24 2165
rect 58 2131 82 2165
rect 0 2097 82 2131
rect 0 2063 24 2097
rect 58 2063 82 2097
rect 0 2029 82 2063
rect 0 1995 24 2029
rect 58 1995 82 2029
rect 0 1961 82 1995
rect 0 1927 24 1961
rect 58 1927 82 1961
rect 0 1893 82 1927
rect 0 1859 24 1893
rect 58 1859 82 1893
rect 0 1825 82 1859
rect 0 1791 24 1825
rect 58 1791 82 1825
rect 0 1757 82 1791
rect 0 1723 24 1757
rect 58 1723 82 1757
rect 0 1689 82 1723
rect 0 1655 24 1689
rect 58 1655 82 1689
rect 0 1621 82 1655
rect 0 1587 24 1621
rect 58 1587 82 1621
rect 0 1553 82 1587
rect 0 1519 24 1553
rect 58 1519 82 1553
rect 0 1485 82 1519
rect 0 1451 24 1485
rect 58 1451 82 1485
rect 0 1417 82 1451
rect 0 1383 24 1417
rect 58 1383 82 1417
rect 0 1349 82 1383
rect 0 1315 24 1349
rect 58 1315 82 1349
rect 0 1281 82 1315
rect 0 1247 24 1281
rect 58 1247 82 1281
rect 0 1213 82 1247
rect 0 1179 24 1213
rect 58 1179 82 1213
rect 0 1145 82 1179
rect 0 1111 24 1145
rect 58 1111 82 1145
rect 0 1077 82 1111
rect 0 1043 24 1077
rect 58 1043 82 1077
rect 0 1009 82 1043
rect 0 975 24 1009
rect 58 975 82 1009
rect 0 941 82 975
rect 0 907 24 941
rect 58 907 82 941
rect 0 873 82 907
rect 0 839 24 873
rect 58 839 82 873
rect 0 805 82 839
rect 0 771 24 805
rect 58 771 82 805
rect 0 737 82 771
rect 0 703 24 737
rect 58 703 82 737
rect 0 669 82 703
rect 0 635 24 669
rect 58 635 82 669
rect 0 601 82 635
rect 0 567 24 601
rect 58 567 82 601
rect 0 533 82 567
rect 0 499 24 533
rect 58 499 82 533
rect 0 465 82 499
rect 0 431 24 465
rect 58 431 82 465
rect 0 397 82 431
rect 0 363 24 397
rect 58 363 82 397
rect 0 329 82 363
rect 0 295 24 329
rect 58 295 82 329
rect 0 261 82 295
rect 0 227 24 261
rect 58 227 82 261
rect 0 193 82 227
rect 0 159 24 193
rect 58 159 82 193
rect 0 125 82 159
rect 0 91 24 125
rect 58 91 82 125
rect 0 57 82 91
rect 0 23 24 57
rect 58 23 82 57
rect 0 0 82 23
<< psubdiffcont >>
rect 24 12943 58 12977
rect 24 12875 58 12909
rect 24 12807 58 12841
rect 24 12739 58 12773
rect 24 12671 58 12705
rect 24 12603 58 12637
rect 24 12535 58 12569
rect 24 12467 58 12501
rect 24 12399 58 12433
rect 24 12331 58 12365
rect 24 12263 58 12297
rect 24 12195 58 12229
rect 24 12127 58 12161
rect 24 12059 58 12093
rect 24 11991 58 12025
rect 24 11923 58 11957
rect 24 11855 58 11889
rect 24 11787 58 11821
rect 24 11719 58 11753
rect 24 11651 58 11685
rect 24 11583 58 11617
rect 24 11515 58 11549
rect 24 11447 58 11481
rect 24 11379 58 11413
rect 24 11311 58 11345
rect 24 11243 58 11277
rect 24 11175 58 11209
rect 24 11107 58 11141
rect 24 11039 58 11073
rect 24 10971 58 11005
rect 24 10903 58 10937
rect 24 10835 58 10869
rect 24 10767 58 10801
rect 24 10699 58 10733
rect 24 10631 58 10665
rect 24 10563 58 10597
rect 24 10495 58 10529
rect 24 10427 58 10461
rect 24 10359 58 10393
rect 24 10291 58 10325
rect 24 10223 58 10257
rect 24 10155 58 10189
rect 24 10087 58 10121
rect 24 10019 58 10053
rect 24 9951 58 9985
rect 24 9883 58 9917
rect 24 9815 58 9849
rect 24 9747 58 9781
rect 24 9679 58 9713
rect 24 9611 58 9645
rect 24 9543 58 9577
rect 24 9475 58 9509
rect 24 9407 58 9441
rect 24 9339 58 9373
rect 24 9271 58 9305
rect 24 9203 58 9237
rect 24 9135 58 9169
rect 24 9067 58 9101
rect 24 8999 58 9033
rect 24 8931 58 8965
rect 24 8863 58 8897
rect 24 8795 58 8829
rect 24 8727 58 8761
rect 24 8659 58 8693
rect 24 8591 58 8625
rect 24 8523 58 8557
rect 24 8455 58 8489
rect 24 8387 58 8421
rect 24 8319 58 8353
rect 24 8251 58 8285
rect 24 8183 58 8217
rect 24 8115 58 8149
rect 24 8047 58 8081
rect 24 7979 58 8013
rect 24 7911 58 7945
rect 24 7843 58 7877
rect 24 7775 58 7809
rect 24 7707 58 7741
rect 24 7639 58 7673
rect 24 7571 58 7605
rect 24 7503 58 7537
rect 24 7435 58 7469
rect 24 7367 58 7401
rect 24 7299 58 7333
rect 24 7231 58 7265
rect 24 7163 58 7197
rect 24 7095 58 7129
rect 24 7027 58 7061
rect 24 6959 58 6993
rect 24 6891 58 6925
rect 24 6823 58 6857
rect 24 6755 58 6789
rect 24 6687 58 6721
rect 24 6619 58 6653
rect 24 6551 58 6585
rect 24 6483 58 6517
rect 24 6415 58 6449
rect 24 6347 58 6381
rect 24 6279 58 6313
rect 24 6211 58 6245
rect 24 6143 58 6177
rect 24 6075 58 6109
rect 24 6007 58 6041
rect 24 5939 58 5973
rect 24 5871 58 5905
rect 24 5803 58 5837
rect 24 5735 58 5769
rect 24 5667 58 5701
rect 24 5599 58 5633
rect 24 5531 58 5565
rect 24 5463 58 5497
rect 24 5395 58 5429
rect 24 5327 58 5361
rect 24 5259 58 5293
rect 24 5191 58 5225
rect 24 5123 58 5157
rect 24 5055 58 5089
rect 24 4987 58 5021
rect 24 4919 58 4953
rect 24 4851 58 4885
rect 24 4783 58 4817
rect 24 4715 58 4749
rect 24 4647 58 4681
rect 24 4579 58 4613
rect 24 4511 58 4545
rect 24 4443 58 4477
rect 24 4375 58 4409
rect 24 4307 58 4341
rect 24 4239 58 4273
rect 24 4171 58 4205
rect 24 4103 58 4137
rect 24 4035 58 4069
rect 24 3967 58 4001
rect 24 3899 58 3933
rect 24 3831 58 3865
rect 24 3763 58 3797
rect 24 3695 58 3729
rect 24 3627 58 3661
rect 24 3559 58 3593
rect 24 3491 58 3525
rect 24 3423 58 3457
rect 24 3355 58 3389
rect 24 3287 58 3321
rect 24 3219 58 3253
rect 24 3151 58 3185
rect 24 3083 58 3117
rect 24 3015 58 3049
rect 24 2947 58 2981
rect 24 2879 58 2913
rect 24 2811 58 2845
rect 24 2743 58 2777
rect 24 2675 58 2709
rect 24 2607 58 2641
rect 24 2539 58 2573
rect 24 2471 58 2505
rect 24 2403 58 2437
rect 24 2335 58 2369
rect 24 2267 58 2301
rect 24 2199 58 2233
rect 24 2131 58 2165
rect 24 2063 58 2097
rect 24 1995 58 2029
rect 24 1927 58 1961
rect 24 1859 58 1893
rect 24 1791 58 1825
rect 24 1723 58 1757
rect 24 1655 58 1689
rect 24 1587 58 1621
rect 24 1519 58 1553
rect 24 1451 58 1485
rect 24 1383 58 1417
rect 24 1315 58 1349
rect 24 1247 58 1281
rect 24 1179 58 1213
rect 24 1111 58 1145
rect 24 1043 58 1077
rect 24 975 58 1009
rect 24 907 58 941
rect 24 839 58 873
rect 24 771 58 805
rect 24 703 58 737
rect 24 635 58 669
rect 24 567 58 601
rect 24 499 58 533
rect 24 431 58 465
rect 24 363 58 397
rect 24 295 58 329
rect 24 227 58 261
rect 24 159 58 193
rect 24 91 58 125
rect 24 23 58 57
<< locali >>
rect 0 12977 82 13000
rect 0 12943 24 12977
rect 58 12943 82 12977
rect 0 12909 82 12943
rect 0 12875 24 12909
rect 58 12875 82 12909
rect 0 12841 82 12875
rect 0 12807 24 12841
rect 58 12807 82 12841
rect 0 12773 82 12807
rect 0 12739 24 12773
rect 58 12739 82 12773
rect 0 12705 82 12739
rect 0 12671 24 12705
rect 58 12671 82 12705
rect 0 12637 82 12671
rect 0 12603 24 12637
rect 58 12603 82 12637
rect 0 12569 82 12603
rect 0 12535 24 12569
rect 58 12535 82 12569
rect 0 12501 82 12535
rect 0 12467 24 12501
rect 58 12467 82 12501
rect 0 12433 82 12467
rect 0 12399 24 12433
rect 58 12399 82 12433
rect 0 12365 82 12399
rect 0 12331 24 12365
rect 58 12331 82 12365
rect 0 12297 82 12331
rect 0 12263 24 12297
rect 58 12263 82 12297
rect 0 12229 82 12263
rect 0 12195 24 12229
rect 58 12195 82 12229
rect 0 12161 82 12195
rect 0 12127 24 12161
rect 58 12127 82 12161
rect 0 12093 82 12127
rect 0 12059 24 12093
rect 58 12059 82 12093
rect 0 12025 82 12059
rect 0 11991 24 12025
rect 58 11991 82 12025
rect 0 11957 82 11991
rect 0 11923 24 11957
rect 58 11923 82 11957
rect 0 11889 82 11923
rect 0 11855 24 11889
rect 58 11855 82 11889
rect 0 11821 82 11855
rect 0 11787 24 11821
rect 58 11787 82 11821
rect 0 11753 82 11787
rect 0 11719 24 11753
rect 58 11719 82 11753
rect 0 11685 82 11719
rect 0 11651 24 11685
rect 58 11651 82 11685
rect 0 11617 82 11651
rect 0 11583 24 11617
rect 58 11583 82 11617
rect 0 11549 82 11583
rect 0 11515 24 11549
rect 58 11515 82 11549
rect 0 11481 82 11515
rect 0 11447 24 11481
rect 58 11447 82 11481
rect 0 11413 82 11447
rect 0 11379 24 11413
rect 58 11379 82 11413
rect 0 11345 82 11379
rect 0 11311 24 11345
rect 58 11311 82 11345
rect 0 11277 82 11311
rect 0 11243 24 11277
rect 58 11243 82 11277
rect 0 11209 82 11243
rect 0 11175 24 11209
rect 58 11175 82 11209
rect 0 11141 82 11175
rect 0 11107 24 11141
rect 58 11107 82 11141
rect 0 11073 82 11107
rect 0 11039 24 11073
rect 58 11039 82 11073
rect 0 11005 82 11039
rect 0 10971 24 11005
rect 58 10971 82 11005
rect 0 10937 82 10971
rect 0 10903 24 10937
rect 58 10903 82 10937
rect 0 10869 82 10903
rect 0 10835 24 10869
rect 58 10835 82 10869
rect 0 10801 82 10835
rect 0 10767 24 10801
rect 58 10767 82 10801
rect 0 10733 82 10767
rect 0 10699 24 10733
rect 58 10699 82 10733
rect 0 10665 82 10699
rect 0 10631 24 10665
rect 58 10631 82 10665
rect 0 10597 82 10631
rect 0 10563 24 10597
rect 58 10563 82 10597
rect 0 10529 82 10563
rect 0 10495 24 10529
rect 58 10495 82 10529
rect 0 10461 82 10495
rect 0 10427 24 10461
rect 58 10427 82 10461
rect 0 10393 82 10427
rect 0 10359 24 10393
rect 58 10359 82 10393
rect 0 10325 82 10359
rect 0 10291 24 10325
rect 58 10291 82 10325
rect 0 10257 82 10291
rect 0 10223 24 10257
rect 58 10223 82 10257
rect 0 10189 82 10223
rect 0 10155 24 10189
rect 58 10155 82 10189
rect 0 10121 82 10155
rect 0 10087 24 10121
rect 58 10087 82 10121
rect 0 10053 82 10087
rect 0 10019 24 10053
rect 58 10019 82 10053
rect 0 9985 82 10019
rect 0 9951 24 9985
rect 58 9951 82 9985
rect 0 9917 82 9951
rect 0 9883 24 9917
rect 58 9883 82 9917
rect 0 9849 82 9883
rect 0 9815 24 9849
rect 58 9815 82 9849
rect 0 9781 82 9815
rect 0 9747 24 9781
rect 58 9747 82 9781
rect 0 9713 82 9747
rect 0 9679 24 9713
rect 58 9679 82 9713
rect 0 9645 82 9679
rect 0 9611 24 9645
rect 58 9611 82 9645
rect 0 9577 82 9611
rect 0 9543 24 9577
rect 58 9543 82 9577
rect 0 9509 82 9543
rect 0 9475 24 9509
rect 58 9475 82 9509
rect 0 9441 82 9475
rect 0 9407 24 9441
rect 58 9407 82 9441
rect 0 9373 82 9407
rect 0 9339 24 9373
rect 58 9339 82 9373
rect 0 9305 82 9339
rect 0 9271 24 9305
rect 58 9271 82 9305
rect 0 9237 82 9271
rect 0 9203 24 9237
rect 58 9203 82 9237
rect 0 9169 82 9203
rect 0 9135 24 9169
rect 58 9135 82 9169
rect 0 9101 82 9135
rect 0 9067 24 9101
rect 58 9067 82 9101
rect 0 9033 82 9067
rect 0 8999 24 9033
rect 58 8999 82 9033
rect 0 8965 82 8999
rect 0 8931 24 8965
rect 58 8931 82 8965
rect 0 8897 82 8931
rect 0 8863 24 8897
rect 58 8863 82 8897
rect 0 8829 82 8863
rect 0 8795 24 8829
rect 58 8795 82 8829
rect 0 8761 82 8795
rect 0 8727 24 8761
rect 58 8727 82 8761
rect 0 8693 82 8727
rect 0 8659 24 8693
rect 58 8659 82 8693
rect 0 8625 82 8659
rect 0 8591 24 8625
rect 58 8591 82 8625
rect 0 8557 82 8591
rect 0 8523 24 8557
rect 58 8523 82 8557
rect 0 8489 82 8523
rect 0 8455 24 8489
rect 58 8455 82 8489
rect 0 8421 82 8455
rect 0 8387 24 8421
rect 58 8387 82 8421
rect 0 8353 82 8387
rect 0 8319 24 8353
rect 58 8319 82 8353
rect 0 8285 82 8319
rect 0 8251 24 8285
rect 58 8251 82 8285
rect 0 8217 82 8251
rect 0 8183 24 8217
rect 58 8183 82 8217
rect 0 8149 82 8183
rect 0 8115 24 8149
rect 58 8115 82 8149
rect 0 8081 82 8115
rect 0 8047 24 8081
rect 58 8047 82 8081
rect 0 8013 82 8047
rect 0 7979 24 8013
rect 58 7979 82 8013
rect 0 7945 82 7979
rect 0 7911 24 7945
rect 58 7911 82 7945
rect 0 7877 82 7911
rect 0 7843 24 7877
rect 58 7843 82 7877
rect 0 7809 82 7843
rect 0 7775 24 7809
rect 58 7775 82 7809
rect 0 7741 82 7775
rect 0 7707 24 7741
rect 58 7707 82 7741
rect 0 7673 82 7707
rect 0 7639 24 7673
rect 58 7639 82 7673
rect 0 7605 82 7639
rect 0 7571 24 7605
rect 58 7571 82 7605
rect 0 7537 82 7571
rect 0 7503 24 7537
rect 58 7503 82 7537
rect 0 7469 82 7503
rect 0 7435 24 7469
rect 58 7435 82 7469
rect 0 7401 82 7435
rect 0 7367 24 7401
rect 58 7367 82 7401
rect 0 7333 82 7367
rect 0 7299 24 7333
rect 58 7299 82 7333
rect 0 7265 82 7299
rect 0 7231 24 7265
rect 58 7231 82 7265
rect 0 7197 82 7231
rect 0 7163 24 7197
rect 58 7163 82 7197
rect 0 7129 82 7163
rect 0 7095 24 7129
rect 58 7095 82 7129
rect 0 7061 82 7095
rect 0 7027 24 7061
rect 58 7027 82 7061
rect 0 6993 82 7027
rect 0 6959 24 6993
rect 58 6959 82 6993
rect 0 6925 82 6959
rect 0 6891 24 6925
rect 58 6891 82 6925
rect 0 6857 82 6891
rect 0 6823 24 6857
rect 58 6823 82 6857
rect 0 6789 82 6823
rect 0 6755 24 6789
rect 58 6755 82 6789
rect 0 6721 82 6755
rect 0 6687 24 6721
rect 58 6687 82 6721
rect 0 6653 82 6687
rect 0 6619 24 6653
rect 58 6619 82 6653
rect 0 6585 82 6619
rect 0 6551 24 6585
rect 58 6551 82 6585
rect 0 6517 82 6551
rect 0 6483 24 6517
rect 58 6483 82 6517
rect 0 6449 82 6483
rect 0 6415 24 6449
rect 58 6415 82 6449
rect 0 6381 82 6415
rect 0 6347 24 6381
rect 58 6347 82 6381
rect 0 6313 82 6347
rect 0 6279 24 6313
rect 58 6279 82 6313
rect 0 6245 82 6279
rect 0 6211 24 6245
rect 58 6211 82 6245
rect 0 6177 82 6211
rect 0 6143 24 6177
rect 58 6143 82 6177
rect 0 6109 82 6143
rect 0 6075 24 6109
rect 58 6075 82 6109
rect 0 6041 82 6075
rect 0 6007 24 6041
rect 58 6007 82 6041
rect 0 5973 82 6007
rect 0 5939 24 5973
rect 58 5939 82 5973
rect 0 5905 82 5939
rect 0 5871 24 5905
rect 58 5871 82 5905
rect 0 5837 82 5871
rect 0 5803 24 5837
rect 58 5803 82 5837
rect 0 5769 82 5803
rect 0 5735 24 5769
rect 58 5735 82 5769
rect 0 5701 82 5735
rect 0 5667 24 5701
rect 58 5667 82 5701
rect 0 5633 82 5667
rect 0 5599 24 5633
rect 58 5599 82 5633
rect 0 5565 82 5599
rect 0 5531 24 5565
rect 58 5531 82 5565
rect 0 5497 82 5531
rect 0 5463 24 5497
rect 58 5463 82 5497
rect 0 5429 82 5463
rect 0 5395 24 5429
rect 58 5395 82 5429
rect 0 5361 82 5395
rect 0 5327 24 5361
rect 58 5327 82 5361
rect 0 5293 82 5327
rect 0 5259 24 5293
rect 58 5259 82 5293
rect 0 5225 82 5259
rect 0 5191 24 5225
rect 58 5191 82 5225
rect 0 5157 82 5191
rect 0 5123 24 5157
rect 58 5123 82 5157
rect 0 5089 82 5123
rect 0 5055 24 5089
rect 58 5055 82 5089
rect 0 5021 82 5055
rect 0 4987 24 5021
rect 58 4987 82 5021
rect 0 4953 82 4987
rect 0 4919 24 4953
rect 58 4919 82 4953
rect 0 4885 82 4919
rect 0 4851 24 4885
rect 58 4851 82 4885
rect 0 4817 82 4851
rect 0 4783 24 4817
rect 58 4783 82 4817
rect 0 4749 82 4783
rect 0 4715 24 4749
rect 58 4715 82 4749
rect 0 4681 82 4715
rect 0 4647 24 4681
rect 58 4647 82 4681
rect 0 4613 82 4647
rect 0 4579 24 4613
rect 58 4579 82 4613
rect 0 4545 82 4579
rect 0 4511 24 4545
rect 58 4511 82 4545
rect 0 4477 82 4511
rect 0 4443 24 4477
rect 58 4443 82 4477
rect 0 4409 82 4443
rect 0 4375 24 4409
rect 58 4375 82 4409
rect 0 4341 82 4375
rect 0 4307 24 4341
rect 58 4307 82 4341
rect 0 4273 82 4307
rect 0 4239 24 4273
rect 58 4239 82 4273
rect 0 4205 82 4239
rect 0 4171 24 4205
rect 58 4171 82 4205
rect 0 4137 82 4171
rect 0 4103 24 4137
rect 58 4103 82 4137
rect 0 4069 82 4103
rect 0 4035 24 4069
rect 58 4035 82 4069
rect 0 4001 82 4035
rect 0 3967 24 4001
rect 58 3967 82 4001
rect 0 3933 82 3967
rect 0 3899 24 3933
rect 58 3899 82 3933
rect 0 3865 82 3899
rect 0 3831 24 3865
rect 58 3831 82 3865
rect 0 3797 82 3831
rect 0 3763 24 3797
rect 58 3763 82 3797
rect 0 3729 82 3763
rect 0 3695 24 3729
rect 58 3695 82 3729
rect 0 3661 82 3695
rect 0 3627 24 3661
rect 58 3627 82 3661
rect 0 3593 82 3627
rect 0 3559 24 3593
rect 58 3559 82 3593
rect 0 3525 82 3559
rect 0 3491 24 3525
rect 58 3491 82 3525
rect 0 3457 82 3491
rect 0 3423 24 3457
rect 58 3423 82 3457
rect 0 3389 82 3423
rect 0 3355 24 3389
rect 58 3355 82 3389
rect 0 3321 82 3355
rect 0 3287 24 3321
rect 58 3287 82 3321
rect 0 3253 82 3287
rect 0 3219 24 3253
rect 58 3219 82 3253
rect 0 3185 82 3219
rect 0 3151 24 3185
rect 58 3151 82 3185
rect 0 3117 82 3151
rect 0 3083 24 3117
rect 58 3083 82 3117
rect 0 3049 82 3083
rect 0 3015 24 3049
rect 58 3015 82 3049
rect 0 2981 82 3015
rect 0 2947 24 2981
rect 58 2947 82 2981
rect 0 2913 82 2947
rect 0 2879 24 2913
rect 58 2879 82 2913
rect 0 2845 82 2879
rect 0 2811 24 2845
rect 58 2811 82 2845
rect 0 2777 82 2811
rect 0 2743 24 2777
rect 58 2743 82 2777
rect 0 2709 82 2743
rect 0 2675 24 2709
rect 58 2675 82 2709
rect 0 2641 82 2675
rect 0 2607 24 2641
rect 58 2607 82 2641
rect 0 2573 82 2607
rect 0 2539 24 2573
rect 58 2539 82 2573
rect 0 2505 82 2539
rect 0 2471 24 2505
rect 58 2471 82 2505
rect 0 2437 82 2471
rect 0 2403 24 2437
rect 58 2403 82 2437
rect 0 2369 82 2403
rect 0 2335 24 2369
rect 58 2335 82 2369
rect 0 2301 82 2335
rect 0 2267 24 2301
rect 58 2267 82 2301
rect 0 2233 82 2267
rect 0 2199 24 2233
rect 58 2199 82 2233
rect 0 2165 82 2199
rect 0 2131 24 2165
rect 58 2131 82 2165
rect 0 2097 82 2131
rect 0 2063 24 2097
rect 58 2063 82 2097
rect 0 2029 82 2063
rect 0 1995 24 2029
rect 58 1995 82 2029
rect 0 1961 82 1995
rect 0 1927 24 1961
rect 58 1927 82 1961
rect 0 1893 82 1927
rect 0 1859 24 1893
rect 58 1859 82 1893
rect 0 1825 82 1859
rect 0 1791 24 1825
rect 58 1791 82 1825
rect 0 1757 82 1791
rect 0 1723 24 1757
rect 58 1723 82 1757
rect 0 1689 82 1723
rect 0 1655 24 1689
rect 58 1655 82 1689
rect 0 1621 82 1655
rect 0 1587 24 1621
rect 58 1587 82 1621
rect 0 1553 82 1587
rect 0 1519 24 1553
rect 58 1519 82 1553
rect 0 1485 82 1519
rect 0 1451 24 1485
rect 58 1451 82 1485
rect 0 1417 82 1451
rect 0 1383 24 1417
rect 58 1383 82 1417
rect 0 1349 82 1383
rect 0 1315 24 1349
rect 58 1315 82 1349
rect 0 1281 82 1315
rect 0 1247 24 1281
rect 58 1247 82 1281
rect 0 1213 82 1247
rect 0 1179 24 1213
rect 58 1179 82 1213
rect 0 1145 82 1179
rect 0 1111 24 1145
rect 58 1111 82 1145
rect 0 1077 82 1111
rect 0 1043 24 1077
rect 58 1043 82 1077
rect 0 1009 82 1043
rect 0 975 24 1009
rect 58 975 82 1009
rect 0 941 82 975
rect 0 907 24 941
rect 58 907 82 941
rect 0 873 82 907
rect 0 839 24 873
rect 58 839 82 873
rect 0 805 82 839
rect 0 771 24 805
rect 58 771 82 805
rect 0 737 82 771
rect 0 703 24 737
rect 58 703 82 737
rect 0 669 82 703
rect 0 635 24 669
rect 58 635 82 669
rect 0 601 82 635
rect 0 567 24 601
rect 58 567 82 601
rect 0 533 82 567
rect 0 499 24 533
rect 58 499 82 533
rect 0 465 82 499
rect 0 431 24 465
rect 58 431 82 465
rect 0 397 82 431
rect 0 363 24 397
rect 58 363 82 397
rect 0 329 82 363
rect 0 295 24 329
rect 58 295 82 329
rect 0 261 82 295
rect 0 227 24 261
rect 58 227 82 261
rect 0 193 82 227
rect 0 159 24 193
rect 58 159 82 193
rect 0 125 82 159
rect 0 91 24 125
rect 58 91 82 125
rect 0 57 82 91
rect 0 23 24 57
rect 58 23 82 57
rect 0 0 82 23
<< end >>
