magic
tech sky130a
timestamp 1739287221
<< checkpaint >>
rect -1070 -221 1054 382
use pfetx241 pfetx241_1
timestamp 1739287221
transform 1 0 -364 0 1 -133
box -47 -88 757 204
use pfetx241 pfetx241_2
timestamp 1739287221
transform 1 0 -363 0 1 178
box -47 -88 757 204
use pfet pfet_1
timestamp 1739287221
transform 1 0 317 0 1 -133
box -47 -88 407 204
use pfet pfet_2
timestamp 1739287221
transform 1 0 317 0 1 178
box -47 -88 407 204
use pfet pfet_3
timestamp 1739287221
transform 1 0 -694 0 1 -133
box -47 -88 407 204
use pfet pfet_4
timestamp 1739287221
transform 1 0 -693 0 1 178
box -47 -88 407 204
use pfet pfet_5
timestamp 1739287221
transform 1 0 -1023 0 1 178
box -47 -88 407 204
use pfet pfet_6
timestamp 1739287221
transform 1 0 -1024 0 1 -133
box -47 -88 407 204
use pfet pfet_7
timestamp 1739287221
transform 1 0 647 0 1 -133
box -47 -88 407 204
use pfet pfet_8
timestamp 1739287221
transform 1 0 647 0 1 178
box -47 -88 407 204
<< end >>
