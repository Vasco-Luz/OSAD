magic
tech sky130A
magscale 1 2
timestamp 1693700175
<< pwell >>
rect -1507 -1027 1507 1027
<< mvnmos >>
rect -1279 -831 -1119 769
rect -1061 -831 -901 769
rect -843 -831 -683 769
rect -625 -831 -465 769
rect -407 -831 -247 769
rect -189 -831 -29 769
rect 29 -831 189 769
rect 247 -831 407 769
rect 465 -831 625 769
rect 683 -831 843 769
rect 901 -831 1061 769
rect 1119 -831 1279 769
<< mvndiff >>
rect -1337 757 -1279 769
rect -1337 -819 -1325 757
rect -1291 -819 -1279 757
rect -1337 -831 -1279 -819
rect -1119 757 -1061 769
rect -1119 -819 -1107 757
rect -1073 -819 -1061 757
rect -1119 -831 -1061 -819
rect -901 757 -843 769
rect -901 -819 -889 757
rect -855 -819 -843 757
rect -901 -831 -843 -819
rect -683 757 -625 769
rect -683 -819 -671 757
rect -637 -819 -625 757
rect -683 -831 -625 -819
rect -465 757 -407 769
rect -465 -819 -453 757
rect -419 -819 -407 757
rect -465 -831 -407 -819
rect -247 757 -189 769
rect -247 -819 -235 757
rect -201 -819 -189 757
rect -247 -831 -189 -819
rect -29 757 29 769
rect -29 -819 -17 757
rect 17 -819 29 757
rect -29 -831 29 -819
rect 189 757 247 769
rect 189 -819 201 757
rect 235 -819 247 757
rect 189 -831 247 -819
rect 407 757 465 769
rect 407 -819 419 757
rect 453 -819 465 757
rect 407 -831 465 -819
rect 625 757 683 769
rect 625 -819 637 757
rect 671 -819 683 757
rect 625 -831 683 -819
rect 843 757 901 769
rect 843 -819 855 757
rect 889 -819 901 757
rect 843 -831 901 -819
rect 1061 757 1119 769
rect 1061 -819 1073 757
rect 1107 -819 1119 757
rect 1061 -831 1119 -819
rect 1279 757 1337 769
rect 1279 -819 1291 757
rect 1325 -819 1337 757
rect 1279 -831 1337 -819
<< mvndiffc >>
rect -1325 -819 -1291 757
rect -1107 -819 -1073 757
rect -889 -819 -855 757
rect -671 -819 -637 757
rect -453 -819 -419 757
rect -235 -819 -201 757
rect -17 -819 17 757
rect 201 -819 235 757
rect 419 -819 453 757
rect 637 -819 671 757
rect 855 -819 889 757
rect 1073 -819 1107 757
rect 1291 -819 1325 757
<< mvpsubdiff >>
rect -1471 979 1471 991
rect -1471 945 -1363 979
rect 1363 945 1471 979
rect -1471 933 1471 945
rect -1471 883 -1413 933
rect -1471 -883 -1459 883
rect -1425 -883 -1413 883
rect 1413 883 1471 933
rect -1471 -933 -1413 -883
rect 1413 -883 1425 883
rect 1459 -883 1471 883
rect 1413 -933 1471 -883
rect -1471 -945 1471 -933
rect -1471 -979 -1363 -945
rect 1363 -979 1471 -945
rect -1471 -991 1471 -979
<< mvpsubdiffcont >>
rect -1363 945 1363 979
rect -1459 -883 -1425 883
rect 1425 -883 1459 883
rect -1363 -979 1363 -945
<< poly >>
rect -1247 841 -1151 857
rect -1247 824 -1231 841
rect -1279 807 -1231 824
rect -1167 824 -1151 841
rect -1029 841 -933 857
rect -1029 824 -1013 841
rect -1167 807 -1119 824
rect -1279 769 -1119 807
rect -1061 807 -1013 824
rect -949 824 -933 841
rect -811 841 -715 857
rect -811 824 -795 841
rect -949 807 -901 824
rect -1061 769 -901 807
rect -843 807 -795 824
rect -731 824 -715 841
rect -593 841 -497 857
rect -593 824 -577 841
rect -731 807 -683 824
rect -843 769 -683 807
rect -625 807 -577 824
rect -513 824 -497 841
rect -375 841 -279 857
rect -375 824 -359 841
rect -513 807 -465 824
rect -625 769 -465 807
rect -407 807 -359 824
rect -295 824 -279 841
rect -157 841 -61 857
rect -157 824 -141 841
rect -295 807 -247 824
rect -407 769 -247 807
rect -189 807 -141 824
rect -77 824 -61 841
rect 61 841 157 857
rect 61 824 77 841
rect -77 807 -29 824
rect -189 769 -29 807
rect 29 807 77 824
rect 141 824 157 841
rect 279 841 375 857
rect 279 824 295 841
rect 141 807 189 824
rect 29 769 189 807
rect 247 807 295 824
rect 359 824 375 841
rect 497 841 593 857
rect 497 824 513 841
rect 359 807 407 824
rect 247 769 407 807
rect 465 807 513 824
rect 577 824 593 841
rect 715 841 811 857
rect 715 824 731 841
rect 577 807 625 824
rect 465 769 625 807
rect 683 807 731 824
rect 795 824 811 841
rect 933 841 1029 857
rect 933 824 949 841
rect 795 807 843 824
rect 683 769 843 807
rect 901 807 949 824
rect 1013 824 1029 841
rect 1151 841 1247 857
rect 1151 824 1167 841
rect 1013 807 1061 824
rect 901 769 1061 807
rect 1119 807 1167 824
rect 1231 824 1247 841
rect 1231 807 1279 824
rect 1119 769 1279 807
rect -1279 -857 -1119 -831
rect -1061 -857 -901 -831
rect -843 -857 -683 -831
rect -625 -857 -465 -831
rect -407 -857 -247 -831
rect -189 -857 -29 -831
rect 29 -857 189 -831
rect 247 -857 407 -831
rect 465 -857 625 -831
rect 683 -857 843 -831
rect 901 -857 1061 -831
rect 1119 -857 1279 -831
<< polycont >>
rect -1231 807 -1167 841
rect -1013 807 -949 841
rect -795 807 -731 841
rect -577 807 -513 841
rect -359 807 -295 841
rect -141 807 -77 841
rect 77 807 141 841
rect 295 807 359 841
rect 513 807 577 841
rect 731 807 795 841
rect 949 807 1013 841
rect 1167 807 1231 841
<< locali >>
rect -1459 945 -1363 979
rect 1363 945 1459 979
rect -1459 883 -1425 945
rect 1425 883 1459 945
rect -1247 807 -1231 841
rect -1167 807 -1151 841
rect -1029 807 -1013 841
rect -949 807 -933 841
rect -811 807 -795 841
rect -731 807 -715 841
rect -593 807 -577 841
rect -513 807 -497 841
rect -375 807 -359 841
rect -295 807 -279 841
rect -157 807 -141 841
rect -77 807 -61 841
rect 61 807 77 841
rect 141 807 157 841
rect 279 807 295 841
rect 359 807 375 841
rect 497 807 513 841
rect 577 807 593 841
rect 715 807 731 841
rect 795 807 811 841
rect 933 807 949 841
rect 1013 807 1029 841
rect 1151 807 1167 841
rect 1231 807 1247 841
rect -1325 757 -1291 773
rect -1325 -835 -1291 -819
rect -1107 757 -1073 773
rect -1107 -835 -1073 -819
rect -889 757 -855 773
rect -889 -835 -855 -819
rect -671 757 -637 773
rect -671 -835 -637 -819
rect -453 757 -419 773
rect -453 -835 -419 -819
rect -235 757 -201 773
rect -235 -835 -201 -819
rect -17 757 17 773
rect -17 -835 17 -819
rect 201 757 235 773
rect 201 -835 235 -819
rect 419 757 453 773
rect 419 -835 453 -819
rect 637 757 671 773
rect 637 -835 671 -819
rect 855 757 889 773
rect 855 -835 889 -819
rect 1073 757 1107 773
rect 1073 -835 1107 -819
rect 1291 757 1325 773
rect 1291 -835 1325 -819
rect -1459 -945 -1425 -883
rect 1425 -945 1459 -883
rect -1459 -979 -1363 -945
rect 1363 -979 1459 -945
<< viali >>
rect -1231 807 -1167 841
rect -1013 807 -949 841
rect -795 807 -731 841
rect -577 807 -513 841
rect -359 807 -295 841
rect -141 807 -77 841
rect 77 807 141 841
rect 295 807 359 841
rect 513 807 577 841
rect 731 807 795 841
rect 949 807 1013 841
rect 1167 807 1231 841
rect -1325 -819 -1291 757
rect -1107 -819 -1073 757
rect -889 -819 -855 757
rect -671 -819 -637 757
rect -453 -819 -419 757
rect -235 -819 -201 757
rect -17 -819 17 757
rect 201 -819 235 757
rect 419 -819 453 757
rect 637 -819 671 757
rect 855 -819 889 757
rect 1073 -819 1107 757
rect 1291 -819 1325 757
<< metal1 >>
rect -1243 841 -1155 847
rect -1243 807 -1231 841
rect -1167 807 -1155 841
rect -1243 801 -1155 807
rect -1025 841 -937 847
rect -1025 807 -1013 841
rect -949 807 -937 841
rect -1025 801 -937 807
rect -807 841 -719 847
rect -807 807 -795 841
rect -731 807 -719 841
rect -807 801 -719 807
rect -589 841 -501 847
rect -589 807 -577 841
rect -513 807 -501 841
rect -589 801 -501 807
rect -371 841 -283 847
rect -371 807 -359 841
rect -295 807 -283 841
rect -371 801 -283 807
rect -153 841 -65 847
rect -153 807 -141 841
rect -77 807 -65 841
rect -153 801 -65 807
rect 65 841 153 847
rect 65 807 77 841
rect 141 807 153 841
rect 65 801 153 807
rect 283 841 371 847
rect 283 807 295 841
rect 359 807 371 841
rect 283 801 371 807
rect 501 841 589 847
rect 501 807 513 841
rect 577 807 589 841
rect 501 801 589 807
rect 719 841 807 847
rect 719 807 731 841
rect 795 807 807 841
rect 719 801 807 807
rect 937 841 1025 847
rect 937 807 949 841
rect 1013 807 1025 841
rect 937 801 1025 807
rect 1155 841 1243 847
rect 1155 807 1167 841
rect 1231 807 1243 841
rect 1155 801 1243 807
rect -1331 757 -1285 769
rect -1331 -819 -1325 757
rect -1291 -819 -1285 757
rect -1331 -831 -1285 -819
rect -1113 757 -1067 769
rect -1113 -819 -1107 757
rect -1073 -819 -1067 757
rect -1113 -831 -1067 -819
rect -895 757 -849 769
rect -895 -819 -889 757
rect -855 -819 -849 757
rect -895 -831 -849 -819
rect -677 757 -631 769
rect -677 -819 -671 757
rect -637 -819 -631 757
rect -677 -831 -631 -819
rect -459 757 -413 769
rect -459 -819 -453 757
rect -419 -819 -413 757
rect -459 -831 -413 -819
rect -241 757 -195 769
rect -241 -819 -235 757
rect -201 -819 -195 757
rect -241 -831 -195 -819
rect -23 757 23 769
rect -23 -819 -17 757
rect 17 -819 23 757
rect -23 -831 23 -819
rect 195 757 241 769
rect 195 -819 201 757
rect 235 -819 241 757
rect 195 -831 241 -819
rect 413 757 459 769
rect 413 -819 419 757
rect 453 -819 459 757
rect 413 -831 459 -819
rect 631 757 677 769
rect 631 -819 637 757
rect 671 -819 677 757
rect 631 -831 677 -819
rect 849 757 895 769
rect 849 -819 855 757
rect 889 -819 895 757
rect 849 -831 895 -819
rect 1067 757 1113 769
rect 1067 -819 1073 757
rect 1107 -819 1113 757
rect 1067 -831 1113 -819
rect 1285 757 1331 769
rect 1285 -819 1291 757
rect 1325 -819 1331 757
rect 1285 -831 1331 -819
<< properties >>
string FIXED_BBOX -1442 -962 1442 962
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 8 l 0.8 m 1 nf 12 diffcov 100 polycov 50 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
