** sch_path: /foss/designs/OSAD/Learning/single_ended_amplifiers/Design_and_Analysis_of_Two-Stage_CMOS_Operational_Amplifier_for_Fluorescence_Signal_Processing_sky130_5V/klayout_layout/Pmos_current_mirror.sch
.subckt Pmos_current_mirror VDD IA IB IC ID
*.PININFO VDD:B IA:B IB:B IC:B ID:B
XM2 IB IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2.2 W='1 * 2 ' nf=2 m=2
XM3 IA IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2.2 W='1 * 2 ' nf=2 m=2
XM4 IC IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2.2 W='1 * 2 ' nf=2 m=8
XM7 ID IA VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2.2 W='1 * 2 ' nf=2 m=16
XM1 IA VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2.2 W='1 * 1 ' nf=1 m=4
XM5 VDD VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2.2 W='1 * 1 ' nf=1 m=4
.ends
.end
