** sch_path: /foss/designs/OSAD/my_ip/testneches_ihp-sg13g2/single_ended_OTAS_testbenches/tb.sch
**.subckt tb
V1 VDD GND 3.3
V2 VSS GND 0
V3 net1 VSS 1.65
V4 VIN+ net1 ac 0.5 sin (0 1m 100k)
V5 VIN- net1 ac -0.5
x1 VDD VSS VIN- VIN+ VOUT amp001_3_3_ihp-sg13g2
C2 VOUT VSS 10p m=1
**** begin user architecture code

.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerHBT.lib hbt_typ


.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerRES.lib res_typ



.param temp=27
.control
op
ac dec 10 1 100G
set appendwrite
write tb.raw
plot db(v(VOUT)) (180*ph(v(VOUT))/pi)
dc V4 0 3.3 0.001
set appendwrite
tran 10ns 50u
set appendwrite
write tb.raw
plot v(VOUT) V(VIN+)


.endc


**** end user architecture code
**.ends

* expanding   symbol:  ihp-sg13g2/Amplifiers/amp001_3_3_ihp-sg13g2.sym # of pins=5
** sym_path: /foss/designs/OSAD/my_ip/LIB/ihp-sg13g2/Amplifiers/amp001_3_3_ihp-sg13g2.sym
** sch_path: /foss/designs/OSAD/my_ip/LIB/ihp-sg13g2/Amplifiers/amp001_3_3_ihp-sg13g2.sch
.subckt amp001_3_3_ihp-sg13g2 VDD VSS VIN- VIN+ VOUT
*.iopin VDD
*.iopin VSS
*.iopin VIN-
*.iopin VIN+
*.iopin VOUT
XQ1 net1 VIN+ net2 VSS npn13G2 Nx=1
XR1 net1 VDD rhigh w=1e-6 l=2e-6 m=1 b=0
XR2 VSS net2 rppd w=0.5e-6 l=1.5e-6 m=1 b=0
XQ2 VDD VIN- net2 VSS npn13G2 Nx=1
XQ6 VOUT net1 net3 pnpMPA a={ 1.0u * 2.0u } p={ ( 1.0u + 2.0u ) * 2 } m=1
XR7 net3 VDD rhigh w=2e-6 l=0.5e-6 m=1 b=0
XR8 VSS VOUT rhigh w=0.5e-6 l=5.4e-6 m=1 b=0
.ends

.GLOBAL GND
.end
