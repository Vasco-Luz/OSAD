* NGSPICE file created from TOP.ext - technology: sky130A

.subckt TOP VDD VSS VIN- VIN+ VOUT
X0 dif_pair_0/IC dif_pair_0/m1_n4845_5624# dif_pair_0/m1_n4845_5624# dif_pair_0/IC sky130_fd_pr__pfet_01v8_lvt ad=0.5 pd=2.5 as=0.6 ps=4.6 w=2 l=0.7
X1 dif_pair_0/IC VIN+ dif_pair_0/II dif_pair_0/IC sky130_fd_pr__pfet_01v8_lvt ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.7
X2 dif_pair_0/IC VIN+ dif_pair_0/II dif_pair_0/IC sky130_fd_pr__pfet_01v8_lvt ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.7
X3 dif_pair_0/m1_n2497_5701# dif_pair_0/m1_n2497_5701# dif_pair_0/IC dif_pair_0/IC sky130_fd_pr__pfet_01v8_lvt ad=0.6 pd=4.6 as=0.5 ps=2.5 w=2 l=0.7
X4 dif_pair_0/IH VIN- dif_pair_0/IC dif_pair_0/IC sky130_fd_pr__pfet_01v8_lvt ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.7
X5 dif_pair_0/IH VIN- dif_pair_0/IC dif_pair_0/IC sky130_fd_pr__pfet_01v8_lvt ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.7
X6 dif_pair_0/II VIN+ dif_pair_0/IC dif_pair_0/IC sky130_fd_pr__pfet_01v8_lvt ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.7
X7 dif_pair_0/IC VIN- dif_pair_0/IH dif_pair_0/IC sky130_fd_pr__pfet_01v8_lvt ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.7
X8 dif_pair_0/IC VIN- dif_pair_0/IH dif_pair_0/IC sky130_fd_pr__pfet_01v8_lvt ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.7
X9 dif_pair_0/II VIN+ dif_pair_0/IC dif_pair_0/IC sky130_fd_pr__pfet_01v8_lvt ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.7
X10 dif_pair_0/IC dif_pair_0/m1_n2497_5948# dif_pair_0/m1_n2497_5948# dif_pair_0/IC sky130_fd_pr__pfet_01v8_lvt ad=14 pd=74 as=0.6 ps=4.6 w=2 l=0.7
X11 dif_pair_0/IC VIN- dif_pair_0/IH dif_pair_0/IC sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=4 ps=20 w=2 l=0.7
X12 dif_pair_0/IC VIN- dif_pair_0/IH dif_pair_0/IC sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2 l=0.7
X13 dif_pair_0/m1_n4845_5948# dif_pair_0/m1_n4845_5948# dif_pair_0/IC dif_pair_0/IC sky130_fd_pr__pfet_01v8_lvt ad=0.6 pd=4.6 as=0 ps=0 w=2 l=0.7
X14 dif_pair_0/II VIN+ dif_pair_0/IC dif_pair_0/IC sky130_fd_pr__pfet_01v8_lvt ad=4 pd=20 as=0 ps=0 w=2 l=0.7
X15 dif_pair_0/II VIN+ dif_pair_0/IC dif_pair_0/IC sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2 l=0.7
X16 dif_pair_0/IH VIN- dif_pair_0/IC dif_pair_0/IC sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2 l=0.7
X17 dif_pair_0/IC VIN+ dif_pair_0/II dif_pair_0/IC sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2 l=0.7
X18 dif_pair_0/IC VIN+ dif_pair_0/II dif_pair_0/IC sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2 l=0.7
X19 dif_pair_0/IH VIN- dif_pair_0/IC dif_pair_0/IC sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2 l=0.7
X20 VSS VSS VSS sky130_fd_pr__res_high_po_0p35 l=2.12
X21 VSS VSS VSS sky130_fd_pr__res_high_po_0p35 l=2.12
X22 VSS m1_1967_n2053# VSS sky130_fd_pr__res_high_po_0p35 l=2.12
X23 m1_1713_n2884# m1_1967_n2053# VSS sky130_fd_pr__res_high_po_0p35 l=2.12
X24 m1_1713_n2884# m1_1459_n2053# VSS sky130_fd_pr__res_high_po_0p35 l=2.12
X25 m1_1205_n2884# m1_1459_n2053# VSS sky130_fd_pr__res_high_po_0p35 l=2.12
X26 m1_1205_n2884# m1_951_n2053# VSS sky130_fd_pr__res_high_po_0p35 l=2.12
X27 m1_697_n2884# m1_951_n2053# VSS sky130_fd_pr__res_high_po_0p35 l=2.12
X28 m1_697_n2884# m1_493_n2053# VSS sky130_fd_pr__res_high_po_0p35 l=2.12
X29 lower_NMOS_0/IG m1_493_n2053# VSS sky130_fd_pr__res_high_po_0p35 l=2.12
X30 lower_NMOS_0/IF lower_NMOS_0/IE lower_NMOS_0/IG VSS sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=4
X31 lower_NMOS_0/IE VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.3 ps=2.6 w=1 l=4
X32 lower_NMOS_0/IF lower_NMOS_0/IE lower_NMOS_0/IG VSS sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=4
X33 lower_NMOS_0/IG lower_NMOS_0/IE lower_NMOS_0/IF VSS sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=4
X34 lower_NMOS_0/IE lower_NMOS_0/IE VSS VSS sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=4
X35 lower_NMOS_0/IG lower_NMOS_0/IE lower_NMOS_0/IF VSS sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=4
X36 VSS lower_NMOS_0/IE lower_NMOS_0/IE VSS sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=4
X37 lower_NMOS_0/IG lower_NMOS_0/IE lower_NMOS_0/IF VSS sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=4
X38 lower_NMOS_0/IG lower_NMOS_0/IE lower_NMOS_0/IF VSS sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=4
X39 lower_NMOS_0/IF VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=4
X40 lower_NMOS_0/IF lower_NMOS_0/IE lower_NMOS_0/IG VSS sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=4
X41 VSS VSS lower_NMOS_0/IF VSS sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=4
X42 VSS VSS lower_NMOS_0/IE VSS sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.25 ps=1.5 w=1 l=4
X43 lower_NMOS_0/IF lower_NMOS_0/IE lower_NMOS_0/IG VSS sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=4
X44 lower_NMOS_0/IF lower_NMOS_0/IE lower_NMOS_0/IG VSS sky130_fd_pr__nfet_01v8 ad=5.5 pd=33 as=4 ps=24 w=1 l=4
X45 lower_NMOS_0/IE VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=4 pd=24 as=13.8 ps=91.4 w=1 l=4
X46 lower_NMOS_0/IF lower_NMOS_0/IE lower_NMOS_0/IG VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=4
X47 lower_NMOS_0/IG lower_NMOS_0/IE lower_NMOS_0/IF VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=4
X48 lower_NMOS_0/IE lower_NMOS_0/IE VSS VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=4
X49 lower_NMOS_0/IG lower_NMOS_0/IE lower_NMOS_0/IF VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=4
X50 VSS lower_NMOS_0/IE lower_NMOS_0/IE VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=4
X51 lower_NMOS_0/IG lower_NMOS_0/IE lower_NMOS_0/IF VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=4
X52 lower_NMOS_0/IG lower_NMOS_0/IE lower_NMOS_0/IF VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=4
X53 lower_NMOS_0/IF VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=4
X54 lower_NMOS_0/IF lower_NMOS_0/IE lower_NMOS_0/IG VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=4
X55 VSS VSS lower_NMOS_0/IF VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=4
X56 VSS VSS lower_NMOS_0/IE VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=4
X57 lower_NMOS_0/IF lower_NMOS_0/IE lower_NMOS_0/IG VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=4
X58 VOUT m1_9568_n4684# sky130_fd_pr__cap_mim_m3_1 l=6.5 w=6.5
X59 VOUT m1_9568_n4684# sky130_fd_pr__cap_mim_m3_1 l=6.5 w=6.5
X60 VOUT m1_9568_n4684# sky130_fd_pr__cap_mim_m3_1 l=6.5 w=6.5
X61 VOUT m1_9568_n4684# sky130_fd_pr__cap_mim_m3_1 l=6.5 w=6.5
X62 dif_pair_0/IH dif_pair_0/IH VSS VSS sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X63 VSS dif_pair_0/IH dif_pair_0/II VSS sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X64 dif_pair_0/IH VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.3 ps=2.6 w=1 l=2
X65 dif_pair_0/II dif_pair_0/IH VSS VSS sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X66 VSS dif_pair_0/IH dif_pair_0/IH VSS sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X67 VSS VSS dif_pair_0/IH VSS sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.25 ps=1.5 w=1 l=2
X68 dif_pair_0/IH dif_pair_0/IH VSS VSS sky130_fd_pr__nfet_01v8 ad=2 pd=12 as=0 ps=0 w=1 l=2
X69 VSS dif_pair_0/IH dif_pair_0/II VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=2.2 ps=15.2 w=1 l=2
X70 dif_pair_0/IH VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=2
X71 dif_pair_0/II dif_pair_0/IH VSS VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=2
X72 VSS dif_pair_0/IH dif_pair_0/IH VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=2
X73 VSS VSS dif_pair_0/IH VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=2
X74 VOUT dif_pair_0/II VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.5
X75 VSS dif_pair_0/II VOUT VSS sky130_fd_pr__nfet_01v8_lvt ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.5
X76 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.5 pd=2.5 as=0.6 ps=4.6 w=2 l=0.5
X77 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.6 pd=4.6 as=0.5 ps=2.5 w=2 l=0.5
X78 VSS dif_pair_0/II VOUT VSS sky130_fd_pr__nfet_01v8_lvt ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.5
X79 VOUT dif_pair_0/II VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.5
X80 VOUT Upper_Nmos_0/IA VDD VDD sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X81 Upper_Nmos_0/IA VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.3 ps=2.6 w=1 l=2
X82 VOUT Upper_Nmos_0/IA VDD VDD sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X83 VDD Upper_Nmos_0/IA VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X84 Upper_Nmos_0/IB Upper_Nmos_0/IA VDD VDD sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X85 VDD Upper_Nmos_0/IA VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X86 VOUT Upper_Nmos_0/IA VDD VDD sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X87 VDD Upper_Nmos_0/IA dif_pair_0/IC VDD sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X88 dif_pair_0/IC Upper_Nmos_0/IA VDD VDD sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X89 VOUT Upper_Nmos_0/IA VDD VDD sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X90 VDD Upper_Nmos_0/IA VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X91 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.6 as=0.25 ps=1.5 w=1 l=2
X92 VDD Upper_Nmos_0/IA VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X93 VOUT Upper_Nmos_0/IA VDD VDD sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X94 VDD Upper_Nmos_0/IA dif_pair_0/IC VDD sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X95 VDD Upper_Nmos_0/IA Upper_Nmos_0/IA VDD sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X96 VOUT Upper_Nmos_0/IA VDD VDD sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X97 VDD Upper_Nmos_0/IA VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X98 VDD Upper_Nmos_0/IA dif_pair_0/IC VDD sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X99 dif_pair_0/IC Upper_Nmos_0/IA VDD VDD sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X100 dif_pair_0/IC Upper_Nmos_0/IA VDD VDD sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X101 VDD Upper_Nmos_0/IA VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X102 VOUT Upper_Nmos_0/IA VDD VDD sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X103 VDD VDD Upper_Nmos_0/IA VDD sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X104 VOUT Upper_Nmos_0/IA VDD VDD sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X105 VDD Upper_Nmos_0/IA dif_pair_0/IC VDD sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X106 Upper_Nmos_0/IA Upper_Nmos_0/IA VDD VDD sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X107 dif_pair_0/IC Upper_Nmos_0/IA VDD VDD sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X108 VDD Upper_Nmos_0/IA VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X109 VDD Upper_Nmos_0/IA Upper_Nmos_0/IB VDD sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X110 VDD Upper_Nmos_0/IA VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X111 VOUT Upper_Nmos_0/IA VDD VDD sky130_fd_pr__pfet_01v8 ad=8 pd=48 as=16.2 ps=100.4 w=1 l=2
X112 Upper_Nmos_0/IA VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2 pd=12 as=0 ps=0 w=1 l=2
X113 VOUT Upper_Nmos_0/IA VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=2
X114 VDD Upper_Nmos_0/IA VOUT VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=2
X115 Upper_Nmos_0/IB Upper_Nmos_0/IA VDD VDD sky130_fd_pr__pfet_01v8 ad=1 pd=6 as=0 ps=0 w=1 l=2
X116 VDD Upper_Nmos_0/IA VOUT VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=2
X117 VOUT Upper_Nmos_0/IA VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=2
X118 VDD Upper_Nmos_0/IA dif_pair_0/IC VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=2
X119 dif_pair_0/IC Upper_Nmos_0/IA VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=2
X120 VOUT Upper_Nmos_0/IA VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=2
X121 VDD Upper_Nmos_0/IA VOUT VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=2
X122 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=2
X123 VDD Upper_Nmos_0/IA VOUT VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=2
X124 VOUT Upper_Nmos_0/IA VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=2
X125 VDD Upper_Nmos_0/IA dif_pair_0/IC VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=2
X126 VDD Upper_Nmos_0/IA Upper_Nmos_0/IA VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=2
X127 VOUT Upper_Nmos_0/IA VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=2
X128 VDD Upper_Nmos_0/IA VOUT VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=2
X129 VDD Upper_Nmos_0/IA dif_pair_0/IC VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=2
X130 dif_pair_0/IC Upper_Nmos_0/IA VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=2
X131 dif_pair_0/IC Upper_Nmos_0/IA VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=2
X132 VDD Upper_Nmos_0/IA VOUT VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=2
X133 VOUT Upper_Nmos_0/IA VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=2
X134 VDD VDD Upper_Nmos_0/IA VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=2
X135 VOUT Upper_Nmos_0/IA VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=2
X136 VDD Upper_Nmos_0/IA dif_pair_0/IC VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=2
X137 Upper_Nmos_0/IA Upper_Nmos_0/IA VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=2
X138 dif_pair_0/IC Upper_Nmos_0/IA VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=2
X139 VDD Upper_Nmos_0/IA VOUT VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=2
X140 VDD Upper_Nmos_0/IA Upper_Nmos_0/IB VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=2
X141 VDD Upper_Nmos_0/IA VOUT VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=2
X142 dif_pair_0/II Upper_Nmos_0/IB m1_9568_n4684# VSS sky130_fd_pr__nfet_01v8 ad=0.6 pd=4.6 as=0.5 ps=2.5 w=2 l=2.2
X143 m1_9568_n4684# Upper_Nmos_0/IB dif_pair_0/II VSS sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.6 ps=4.6 w=2 l=2.2
X144 Upper_Nmos_0/IA VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X145 Upper_Nmos_0/IB VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.25 pd=1.5 as=0.3 ps=2.6 w=1 l=2
X146 VSS VSS lower_NMOS_0/IE VSS sky130_fd_pr__nfet_01v8_lvt ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X147 VSS VSS Upper_Nmos_0/IB VSS sky130_fd_pr__nfet_01v8_lvt ad=0.3 pd=2.6 as=0.25 ps=1.5 w=1 l=2
X148 Upper_Nmos_0/IB Upper_Nmos_0/IB lower_NMOS_0/IE VSS sky130_fd_pr__nfet_01v8_lvt ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X149 lower_NMOS_0/IE VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X150 lower_NMOS_0/IE Upper_Nmos_0/IB Upper_Nmos_0/IB VSS sky130_fd_pr__nfet_01v8_lvt ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X151 VSS VSS Upper_Nmos_0/IA VSS sky130_fd_pr__nfet_01v8_lvt ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X152 Upper_Nmos_0/IA Upper_Nmos_0/IB Upper_Nmos_0/nfet_0/a_2460_0# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X153 Upper_Nmos_0/nfet_0/a_2460_0# Upper_Nmos_0/IB Upper_Nmos_0/IA VSS sky130_fd_pr__nfet_01v8_lvt ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=2
X154 Upper_Nmos_0/IA VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=2 pd=12 as=0 ps=0 w=1 l=2
X155 Upper_Nmos_0/IB VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=2 pd=12 as=0 ps=0 w=1 l=2
X156 VSS VSS lower_NMOS_0/IE VSS sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1 l=2
X157 VSS VSS Upper_Nmos_0/IB VSS sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1 l=2
X158 Upper_Nmos_0/IB Upper_Nmos_0/IB lower_NMOS_0/IE VSS sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1 l=2
X159 lower_NMOS_0/IE VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1 l=2
X160 lower_NMOS_0/IE Upper_Nmos_0/IB Upper_Nmos_0/IB VSS sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1 l=2
X161 VSS VSS Upper_Nmos_0/IA VSS sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1 l=2
X162 Upper_Nmos_0/IA Upper_Nmos_0/IB lower_NMOS_0/IF VSS sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1 l=2
X163 lower_NMOS_0/IF Upper_Nmos_0/IB Upper_Nmos_0/IA VSS sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1 l=2
C0 dif_pair_0/IH dif_pair_0/IC 2.56783f
C1 Upper_Nmos_0/IA VOUT 3.61544f
C2 Upper_Nmos_0/IA Upper_Nmos_0/IB 2.58035f
C3 VIN+ VIN- 2.74653f
C4 lower_NMOS_0/IF lower_NMOS_0/IE 6.29946f
C5 VOUT dif_pair_0/IC 5.32644f
C6 VDD Upper_Nmos_0/IA 37.30863f
C7 VSS lower_NMOS_0/IE 10.40228f
C8 VSS m1_9568_n4684# 2.97159f
C9 VDD dif_pair_0/IC 2.53356f
C10 VSS dif_pair_0/IH 2.72891f
C11 m1_9568_n4684# VOUT 19.1651f
C12 dif_pair_0/II dif_pair_0/IC 2.15402f
C13 Upper_Nmos_0/IA dif_pair_0/IC 2.79614f
C14 VSS VOUT 2.98876f
C15 VSS Upper_Nmos_0/IB 5.78101f
C16 dif_pair_0/IH Upper_Nmos_0/IB 2.0653f
C17 lower_NMOS_0/IG lower_NMOS_0/IE 2.42788f
C18 Upper_Nmos_0/IB VOUT 3.94645f
C19 lower_NMOS_0/IF lower_NMOS_0/IG 3.40712f
C20 dif_pair_0/II dif_pair_0/IH 3.23565f
C21 VIN+ dif_pair_0/IC 2.49173f
C22 VIN- dif_pair_0/IC 2.4612f
C23 VDD VOUT 2.67062f
C24 Upper_Nmos_0/IB 0 11.38539f
C25 VOUT 0 6.84386f
C26 Upper_Nmos_0/IA 0 17.23009f
C27 VDD 0 76.51212f
C28 dif_pair_0/IH 0 6.59843f
C29 m1_9568_n4684# 0 6.87714f $ **FLOATING
C30 VSS 0 20.33185f
C31 lower_NMOS_0/IE 0 30.1416f
C32 dif_pair_0/II 0 3.37007f
C33 dif_pair_0/IC 0 16.08201f
.ends
