magic
tech sky130A
magscale 1 2
timestamp 1693699723
<< nwell >>
rect -1537 -662 1537 662
<< mvpmos >>
rect -1279 -436 -1119 364
rect -1061 -436 -901 364
rect -843 -436 -683 364
rect -625 -436 -465 364
rect -407 -436 -247 364
rect -189 -436 -29 364
rect 29 -436 189 364
rect 247 -436 407 364
rect 465 -436 625 364
rect 683 -436 843 364
rect 901 -436 1061 364
rect 1119 -436 1279 364
<< mvpdiff >>
rect -1337 352 -1279 364
rect -1337 -424 -1325 352
rect -1291 -424 -1279 352
rect -1337 -436 -1279 -424
rect -1119 352 -1061 364
rect -1119 -424 -1107 352
rect -1073 -424 -1061 352
rect -1119 -436 -1061 -424
rect -901 352 -843 364
rect -901 -424 -889 352
rect -855 -424 -843 352
rect -901 -436 -843 -424
rect -683 352 -625 364
rect -683 -424 -671 352
rect -637 -424 -625 352
rect -683 -436 -625 -424
rect -465 352 -407 364
rect -465 -424 -453 352
rect -419 -424 -407 352
rect -465 -436 -407 -424
rect -247 352 -189 364
rect -247 -424 -235 352
rect -201 -424 -189 352
rect -247 -436 -189 -424
rect -29 352 29 364
rect -29 -424 -17 352
rect 17 -424 29 352
rect -29 -436 29 -424
rect 189 352 247 364
rect 189 -424 201 352
rect 235 -424 247 352
rect 189 -436 247 -424
rect 407 352 465 364
rect 407 -424 419 352
rect 453 -424 465 352
rect 407 -436 465 -424
rect 625 352 683 364
rect 625 -424 637 352
rect 671 -424 683 352
rect 625 -436 683 -424
rect 843 352 901 364
rect 843 -424 855 352
rect 889 -424 901 352
rect 843 -436 901 -424
rect 1061 352 1119 364
rect 1061 -424 1073 352
rect 1107 -424 1119 352
rect 1061 -436 1119 -424
rect 1279 352 1337 364
rect 1279 -424 1291 352
rect 1325 -424 1337 352
rect 1279 -436 1337 -424
<< mvpdiffc >>
rect -1325 -424 -1291 352
rect -1107 -424 -1073 352
rect -889 -424 -855 352
rect -671 -424 -637 352
rect -453 -424 -419 352
rect -235 -424 -201 352
rect -17 -424 17 352
rect 201 -424 235 352
rect 419 -424 453 352
rect 637 -424 671 352
rect 855 -424 889 352
rect 1073 -424 1107 352
rect 1291 -424 1325 352
<< mvnsubdiff >>
rect -1471 584 1471 596
rect -1471 550 -1363 584
rect 1363 550 1471 584
rect -1471 538 1471 550
rect -1471 488 -1413 538
rect -1471 -488 -1459 488
rect -1425 -488 -1413 488
rect 1413 488 1471 538
rect -1471 -538 -1413 -488
rect 1413 -488 1425 488
rect 1459 -488 1471 488
rect 1413 -538 1471 -488
rect -1471 -550 1471 -538
rect -1471 -584 -1363 -550
rect 1363 -584 1471 -550
rect -1471 -596 1471 -584
<< mvnsubdiffcont >>
rect -1363 550 1363 584
rect -1459 -488 -1425 488
rect 1425 -488 1459 488
rect -1363 -584 1363 -550
<< poly >>
rect -1253 445 -1145 461
rect -1253 428 -1237 445
rect -1279 411 -1237 428
rect -1161 428 -1145 445
rect -1035 445 -927 461
rect -1035 428 -1019 445
rect -1161 411 -1119 428
rect -1279 364 -1119 411
rect -1061 411 -1019 428
rect -943 428 -927 445
rect -817 445 -709 461
rect -817 428 -801 445
rect -943 411 -901 428
rect -1061 364 -901 411
rect -843 411 -801 428
rect -725 428 -709 445
rect -599 445 -491 461
rect -599 428 -583 445
rect -725 411 -683 428
rect -843 364 -683 411
rect -625 411 -583 428
rect -507 428 -491 445
rect -381 445 -273 461
rect -381 428 -365 445
rect -507 411 -465 428
rect -625 364 -465 411
rect -407 411 -365 428
rect -289 428 -273 445
rect -163 445 -55 461
rect -163 428 -147 445
rect -289 411 -247 428
rect -407 364 -247 411
rect -189 411 -147 428
rect -71 428 -55 445
rect 55 445 163 461
rect 55 428 71 445
rect -71 411 -29 428
rect -189 364 -29 411
rect 29 411 71 428
rect 147 428 163 445
rect 273 445 381 461
rect 273 428 289 445
rect 147 411 189 428
rect 29 364 189 411
rect 247 411 289 428
rect 365 428 381 445
rect 491 445 599 461
rect 491 428 507 445
rect 365 411 407 428
rect 247 364 407 411
rect 465 411 507 428
rect 583 428 599 445
rect 709 445 817 461
rect 709 428 725 445
rect 583 411 625 428
rect 465 364 625 411
rect 683 411 725 428
rect 801 428 817 445
rect 927 445 1035 461
rect 927 428 943 445
rect 801 411 843 428
rect 683 364 843 411
rect 901 411 943 428
rect 1019 428 1035 445
rect 1145 445 1253 461
rect 1145 428 1161 445
rect 1019 411 1061 428
rect 901 364 1061 411
rect 1119 411 1161 428
rect 1237 428 1253 445
rect 1237 411 1279 428
rect 1119 364 1279 411
rect -1279 -462 -1119 -436
rect -1061 -462 -901 -436
rect -843 -462 -683 -436
rect -625 -462 -465 -436
rect -407 -462 -247 -436
rect -189 -462 -29 -436
rect 29 -462 189 -436
rect 247 -462 407 -436
rect 465 -462 625 -436
rect 683 -462 843 -436
rect 901 -462 1061 -436
rect 1119 -462 1279 -436
<< polycont >>
rect -1237 411 -1161 445
rect -1019 411 -943 445
rect -801 411 -725 445
rect -583 411 -507 445
rect -365 411 -289 445
rect -147 411 -71 445
rect 71 411 147 445
rect 289 411 365 445
rect 507 411 583 445
rect 725 411 801 445
rect 943 411 1019 445
rect 1161 411 1237 445
<< locali >>
rect -1459 550 -1363 584
rect 1363 550 1459 584
rect -1459 488 -1425 550
rect 1425 488 1459 550
rect -1253 411 -1237 445
rect -1161 411 -1145 445
rect -1035 411 -1019 445
rect -943 411 -927 445
rect -817 411 -801 445
rect -725 411 -709 445
rect -599 411 -583 445
rect -507 411 -491 445
rect -381 411 -365 445
rect -289 411 -273 445
rect -163 411 -147 445
rect -71 411 -55 445
rect 55 411 71 445
rect 147 411 163 445
rect 273 411 289 445
rect 365 411 381 445
rect 491 411 507 445
rect 583 411 599 445
rect 709 411 725 445
rect 801 411 817 445
rect 927 411 943 445
rect 1019 411 1035 445
rect 1145 411 1161 445
rect 1237 411 1253 445
rect -1325 352 -1291 368
rect -1325 -440 -1291 -424
rect -1107 352 -1073 368
rect -1107 -440 -1073 -424
rect -889 352 -855 368
rect -889 -440 -855 -424
rect -671 352 -637 368
rect -671 -440 -637 -424
rect -453 352 -419 368
rect -453 -440 -419 -424
rect -235 352 -201 368
rect -235 -440 -201 -424
rect -17 352 17 368
rect -17 -440 17 -424
rect 201 352 235 368
rect 201 -440 235 -424
rect 419 352 453 368
rect 419 -440 453 -424
rect 637 352 671 368
rect 637 -440 671 -424
rect 855 352 889 368
rect 855 -440 889 -424
rect 1073 352 1107 368
rect 1073 -440 1107 -424
rect 1291 352 1325 368
rect 1291 -440 1325 -424
rect -1459 -550 -1425 -488
rect 1425 -550 1459 -488
rect -1459 -584 -1363 -550
rect 1363 -584 1459 -550
<< viali >>
rect -1237 411 -1161 445
rect -1019 411 -943 445
rect -801 411 -725 445
rect -583 411 -507 445
rect -365 411 -289 445
rect -147 411 -71 445
rect 71 411 147 445
rect 289 411 365 445
rect 507 411 583 445
rect 725 411 801 445
rect 943 411 1019 445
rect 1161 411 1237 445
rect -1325 -424 -1291 352
rect -1107 -424 -1073 352
rect -889 -424 -855 352
rect -671 -424 -637 352
rect -453 -424 -419 352
rect -235 -424 -201 352
rect -17 -424 17 352
rect 201 -424 235 352
rect 419 -424 453 352
rect 637 -424 671 352
rect 855 -424 889 352
rect 1073 -424 1107 352
rect 1291 -424 1325 352
<< metal1 >>
rect -1249 445 -1149 451
rect -1249 411 -1237 445
rect -1161 411 -1149 445
rect -1249 405 -1149 411
rect -1031 445 -931 451
rect -1031 411 -1019 445
rect -943 411 -931 445
rect -1031 405 -931 411
rect -813 445 -713 451
rect -813 411 -801 445
rect -725 411 -713 445
rect -813 405 -713 411
rect -595 445 -495 451
rect -595 411 -583 445
rect -507 411 -495 445
rect -595 405 -495 411
rect -377 445 -277 451
rect -377 411 -365 445
rect -289 411 -277 445
rect -377 405 -277 411
rect -159 445 -59 451
rect -159 411 -147 445
rect -71 411 -59 445
rect -159 405 -59 411
rect 59 445 159 451
rect 59 411 71 445
rect 147 411 159 445
rect 59 405 159 411
rect 277 445 377 451
rect 277 411 289 445
rect 365 411 377 445
rect 277 405 377 411
rect 495 445 595 451
rect 495 411 507 445
rect 583 411 595 445
rect 495 405 595 411
rect 713 445 813 451
rect 713 411 725 445
rect 801 411 813 445
rect 713 405 813 411
rect 931 445 1031 451
rect 931 411 943 445
rect 1019 411 1031 445
rect 931 405 1031 411
rect 1149 445 1249 451
rect 1149 411 1161 445
rect 1237 411 1249 445
rect 1149 405 1249 411
rect -1331 352 -1285 364
rect -1331 -424 -1325 352
rect -1291 -424 -1285 352
rect -1331 -436 -1285 -424
rect -1113 352 -1067 364
rect -1113 -424 -1107 352
rect -1073 -424 -1067 352
rect -1113 -436 -1067 -424
rect -895 352 -849 364
rect -895 -424 -889 352
rect -855 -424 -849 352
rect -895 -436 -849 -424
rect -677 352 -631 364
rect -677 -424 -671 352
rect -637 -424 -631 352
rect -677 -436 -631 -424
rect -459 352 -413 364
rect -459 -424 -453 352
rect -419 -424 -413 352
rect -459 -436 -413 -424
rect -241 352 -195 364
rect -241 -424 -235 352
rect -201 -424 -195 352
rect -241 -436 -195 -424
rect -23 352 23 364
rect -23 -424 -17 352
rect 17 -424 23 352
rect -23 -436 23 -424
rect 195 352 241 364
rect 195 -424 201 352
rect 235 -424 241 352
rect 195 -436 241 -424
rect 413 352 459 364
rect 413 -424 419 352
rect 453 -424 459 352
rect 413 -436 459 -424
rect 631 352 677 364
rect 631 -424 637 352
rect 671 -424 677 352
rect 631 -436 677 -424
rect 849 352 895 364
rect 849 -424 855 352
rect 889 -424 895 352
rect 849 -436 895 -424
rect 1067 352 1113 364
rect 1067 -424 1073 352
rect 1107 -424 1113 352
rect 1067 -436 1113 -424
rect 1285 352 1331 364
rect 1285 -424 1291 352
rect 1325 -424 1331 352
rect 1285 -436 1331 -424
<< properties >>
string FIXED_BBOX -1442 -567 1442 567
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 4 l 0.8 m 1 nf 12 diffcov 100 polycov 60 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 60 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
