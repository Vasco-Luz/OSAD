** sch_path: /home/vasco/Desktop/sky130A/amplifiers/differencial_stage_amps/stange
*+ stages/basic_NMOS_resistive_stage/diferential_stage.sch
**.subckt diferential_stage
XM5 VOUT+ VIN net1 GND sky130_fd_pr__nfet_g5v0d10v5 L=0.7 W=25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 VOUT- VB net1 GND sky130_fd_pr__nfet_g5v0d10v5 L=0.7 W=25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
V1 VDD GND 5
.save i(v1)
V2 VIN GND 2.5
.save i(v2)
V6 VB GND 2.5
.save i(v6)
XM2 net3 net2 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=100 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
Vmeas net1 net3 0
.save i(vmeas)
R5 VOUT+_tran GND 10G m=1
R2 VIN net4 10G m=1
V4 VIN_tran GND ac 1.0 sin (0 100u 100k)
.save i(v4)
C1 VIN_tran net4 1 m=1
R3 VIN net5 10G m=1
C3 net6 net5 1 m=1
V5 net6 GND ac 1.0 sin (0 100u 100k)
.save i(v5)
R4 VOUT+_ac GND 10G m=1
V7 net7 VDD ac 1.0 sin (0 0u 100k)
.save i(v7)
R7 VOUT+_a+ GND 10G m=1
V8 net8 GND ac 1.0 sin (0 0u 100k)
.save i(v8)
R8 VOUT+_a- GND 10G m=1
R9 VB net9 10G m=1
C4 net10 net9 1 m=1
V10 net10 GND ac 1.0 sin (0 100u 100k)
.save i(v10)
XM3 net2 net2 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=100 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
I0 VDD net2 0.2m
XM9 VOUT+ VOUT+ VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 VOUT- VOUT- VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XR6 VOUT+ VOUT- VDD sky130_fd_pr__res_high_po_0p35 L=1*30 mult=1 m=1
x1 VDD GND net4 VB VOUT+_tran differential_stage
x2 VDD GND net5 VB VOUT+_ac differential_stage
x3 net7 GND VIN VB VOUT+_a+ differential_stage
x4 VDD net8 VIN VB VOUT+_a- differential_stage
x5 VDD GND net9 net9 VOUT+_CA differential_stage
**** begin user architecture code

**************************************************************
**************************************************************
**************************************************************
**************************************************************
**************************************************************
*LIBs*********************************************************
**************************************************************
**************************************************************
**************************************************************
**************************************************************
**************************************************************
*.lib /home/vasco/Desktop/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
* chose the corners in the corner file
* tt_mm for mismatch
* ss ff sf fs standart corners
* ll hh lh hl capacitor and resistors corners
* mc for total process variation including corners
**************************************************************
**************************************************************
**************************************************************
**************************************************************
**************************************************************
*Corners/montecarlo options***********************************
**************************************************************
**************************************************************
**************************************************************
**************************************************************
**************************************************************
.TEMP 27
**************************************************************
**************************************************************
**************************************************************
**************************************************************
*SIMULATION and Plots*****************************************
**************************************************************
**************************************************************
**************************************************************
**************************************************************
.control
save all
dc V2 0 5 0.01
*dc simulation
plot v(VOUT-) v(VIN) deriv(v(VOUT-)) v(VOUT+) deriv(v(VOUT+))
*ploting VIN VOUT and the voltage gain
plot i(Vmeas)
*ploting the current for curiosity
tran 1ns 20u
*transient simulation
plot (v(VOUT+_tran))
*simple plot to exemplify the gain
fft v(VOUT+_tran) v(VIN_tran)
*fast fourier transfor
plot mag(v(VOUT+_tran)) mag(v(VIN_tran))
ac dec 20 1 1000G
*simple ac simulation
plot db(v(VOUT+_ac))
plot db(v(VOUT+_a+))
plot db(v(VOUT+_a-))
plot db(v(VOUT+_CA))
plot db((v(VOUT+_ac))/(v(VOUT+_CA)))
plot db((v(VOUT+_ac))/(v(VOUT+_a+)))
plot db((v(VOUT+_ac))/(v(VOUT+_a-)))
.endc


.param mc_mm_switch=0
.param mc_pr_switch=0
.include /home/vasco/Desktop/pdk/sky130A/libs.tech/ngspice/corners/tt.spice
.include /home/vasco/Desktop/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/vasco/Desktop/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/vasco/Desktop/pdk/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends

* expanding   symbol:  /home/vasco/Desktop/sky130A/amplifiers/differencial_stage_amps/stange
*+ stages/basic_NMOS_resistive_stage/differential_stage.sym # of pins=5
** sym_path: /home/vasco/Desktop/sky130A/amplifiers/differencial_stage_amps/stange
*+ stages/basic_NMOS_resistive_stage/differential_stage.sym
** sch_path: /home/vasco/Desktop/sky130A/amplifiers/differencial_stage_amps/stange
*+ stages/basic_NMOS_resistive_stage/differential_stage.sch
.subckt differential_stage VDD VSS VIN+ VIN- VOUT+
*.iopin VDD
*.iopin VSS
*.iopin VIN+
*.iopin VIN-
*.iopin VOUT+
XM5 VOUT+ VIN+ net1 VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.7 W=25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 VOUT- VIN- net1 VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.7 W=25 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 net1 net2 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=100 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 net2 net2 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=100 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
I0 VDD net2 200u
XM9 VOUT+ VOUT+ VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 VOUT- VOUT- VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XR6 VOUT+ VOUT- VDD sky130_fd_pr__res_high_po_0p35 L=1*30 mult=1 m=1
.ends

.GLOBAL GND
.end
