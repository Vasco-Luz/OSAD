magic
tech sky130A
magscale 1 2
timestamp 1740346228
<< error_p >>
rect -324 198 324 202
rect -324 -130 -294 198
rect -258 132 258 136
rect -258 -64 -228 132
rect 228 -64 258 132
rect 294 -130 324 198
<< nwell >>
rect -294 -164 294 198
<< mvpmos >>
rect -200 -64 200 136
<< mvpdiff >>
rect -258 124 -200 136
rect -258 -52 -246 124
rect -212 -52 -200 124
rect -258 -64 -200 -52
rect 200 124 258 136
rect 200 -52 212 124
rect 246 -52 258 124
rect 200 -64 258 -52
<< mvpdiffc >>
rect -246 -52 -212 124
rect 212 -52 246 124
<< poly >>
rect -200 136 200 162
rect -200 -111 200 -64
rect -200 -128 -147 -111
rect -163 -145 -147 -128
rect 147 -128 200 -111
rect 147 -145 163 -128
rect -163 -161 163 -145
<< polycont >>
rect -147 -145 147 -111
<< locali >>
rect -246 124 -212 140
rect -246 -68 -212 -52
rect 212 124 246 140
rect 212 -68 246 -52
rect -164 -111 164 -110
rect -164 -145 -147 -111
rect 147 -145 164 -111
rect -164 -180 164 -145
rect -246 -194 266 -180
rect -246 -228 -234 -194
rect -200 -228 -148 -194
rect -114 -228 266 -194
rect -246 -240 266 -228
<< viali >>
rect -246 -52 -212 124
rect 212 -52 246 124
rect -147 -145 147 -111
rect -234 -228 -200 -194
rect -148 -228 -114 -194
<< metal1 >>
rect 212 136 246 206
rect -252 124 -206 136
rect -252 -52 -246 124
rect -212 -52 -206 124
rect -252 -64 -206 -52
rect 206 124 252 136
rect 206 -52 212 124
rect 246 -52 252 124
rect 206 -64 252 -52
rect -246 -180 -212 -64
rect -159 -111 159 -105
rect -159 -145 -147 -111
rect 147 -145 159 -111
rect -159 -151 159 -145
rect -246 -194 -102 -180
rect -246 -228 -234 -194
rect -200 -228 -148 -194
rect -114 -228 -102 -194
rect -246 -240 -102 -228
<< labels >>
flabel mvpmos -92 -8 82 54 0 FreeSans 800 0 0 0 M3
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1 l 2 m 1 nf 1 diffcov 100 polycov 80 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 80 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
