magic
tech gf180mcuD
magscale 1 10
timestamp 1714262332
<< nwell >>
rect -550 -1358 550 1358
<< pmos >>
rect -300 748 300 1148
rect -300 116 300 516
rect -300 -516 300 -116
rect -300 -1148 300 -748
<< pdiff >>
rect -388 1135 -300 1148
rect -388 761 -375 1135
rect -329 761 -300 1135
rect -388 748 -300 761
rect 300 1135 388 1148
rect 300 761 329 1135
rect 375 761 388 1135
rect 300 748 388 761
rect -388 503 -300 516
rect -388 129 -375 503
rect -329 129 -300 503
rect -388 116 -300 129
rect 300 503 388 516
rect 300 129 329 503
rect 375 129 388 503
rect 300 116 388 129
rect -388 -129 -300 -116
rect -388 -503 -375 -129
rect -329 -503 -300 -129
rect -388 -516 -300 -503
rect 300 -129 388 -116
rect 300 -503 329 -129
rect 375 -503 388 -129
rect 300 -516 388 -503
rect -388 -761 -300 -748
rect -388 -1135 -375 -761
rect -329 -1135 -300 -761
rect -388 -1148 -300 -1135
rect 300 -761 388 -748
rect 300 -1135 329 -761
rect 375 -1135 388 -761
rect 300 -1148 388 -1135
<< pdiffc >>
rect -375 761 -329 1135
rect 329 761 375 1135
rect -375 129 -329 503
rect 329 129 375 503
rect -375 -503 -329 -129
rect 329 -503 375 -129
rect -375 -1135 -329 -761
rect 329 -1135 375 -761
<< nsubdiff >>
rect -526 1262 526 1334
rect -526 1218 -454 1262
rect -526 -1218 -513 1218
rect -467 -1218 -454 1218
rect 454 1218 526 1262
rect -526 -1262 -454 -1218
rect 454 -1218 467 1218
rect 513 -1218 526 1218
rect 454 -1262 526 -1218
rect -526 -1334 526 -1262
<< nsubdiffcont >>
rect -513 -1218 -467 1218
rect 467 -1218 513 1218
<< polysilicon >>
rect -300 1227 300 1240
rect -300 1181 -287 1227
rect 287 1181 300 1227
rect -300 1148 300 1181
rect -300 715 300 748
rect -300 669 -287 715
rect 287 669 300 715
rect -300 656 300 669
rect -300 595 300 608
rect -300 549 -287 595
rect 287 549 300 595
rect -300 516 300 549
rect -300 83 300 116
rect -300 37 -287 83
rect 287 37 300 83
rect -300 24 300 37
rect -300 -37 300 -24
rect -300 -83 -287 -37
rect 287 -83 300 -37
rect -300 -116 300 -83
rect -300 -549 300 -516
rect -300 -595 -287 -549
rect 287 -595 300 -549
rect -300 -608 300 -595
rect -300 -669 300 -656
rect -300 -715 -287 -669
rect 287 -715 300 -669
rect -300 -748 300 -715
rect -300 -1181 300 -1148
rect -300 -1227 -287 -1181
rect 287 -1227 300 -1181
rect -300 -1240 300 -1227
<< polycontact >>
rect -287 1181 287 1227
rect -287 669 287 715
rect -287 549 287 595
rect -287 37 287 83
rect -287 -83 287 -37
rect -287 -595 287 -549
rect -287 -715 287 -669
rect -287 -1227 287 -1181
<< metal1 >>
rect -513 1275 513 1321
rect -513 1218 -467 1275
rect -298 1181 -287 1227
rect 287 1181 298 1227
rect 467 1218 513 1275
rect -375 1135 -329 1146
rect -375 750 -329 761
rect 329 1135 375 1146
rect 329 750 375 761
rect -298 669 -287 715
rect 287 669 298 715
rect -298 549 -287 595
rect 287 549 298 595
rect -375 503 -329 514
rect -375 118 -329 129
rect 329 503 375 514
rect 329 118 375 129
rect -298 37 -287 83
rect 287 37 298 83
rect -298 -83 -287 -37
rect 287 -83 298 -37
rect -375 -129 -329 -118
rect -375 -514 -329 -503
rect 329 -129 375 -118
rect 329 -514 375 -503
rect -298 -595 -287 -549
rect 287 -595 298 -549
rect -298 -715 -287 -669
rect 287 -715 298 -669
rect -375 -761 -329 -750
rect -375 -1146 -329 -1135
rect 329 -761 375 -750
rect 329 -1146 375 -1135
rect -513 -1275 -467 -1218
rect -298 -1227 -287 -1181
rect 287 -1227 298 -1181
rect 467 -1275 513 -1218
rect -513 -1321 513 -1275
<< properties >>
string FIXED_BBOX -490 -1298 490 1298
string gencell pfet_03v3
string library gf180mcu
string parameters w 2.0 l 3.0 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 1 compatible {pfet_03v3 pfet_06v0}
<< end >>
