** sch_path: /foss/designs/OSAD/Learning/fully_differencial/Indirect_Compensation_Techniques_for_Three_Stage_Fully_Differential_Op_amps_IHP130/testbenches/transimpedance_cell_tb_.sch
**.subckt transimpedance_cell_tb_
V1 VDD GND VDD
V2 VSS GND VSS
XM1 net3 net1 VDD VDD sg13_hv_pmos w=1.5u l=3u ng=2 m=2
XM2 net1 net1 VDD VDD sg13_hv_pmos w=1.5u l=3u ng=2 m=2
XM6 net2 VSS VSS VSS sg13_hv_nmos w=4.5u l=2u ng=2 m=2
Vmeas2 VDD net2 0
.save i(vmeas2)
Vmeas1 net3 net4 0
.save i(vmeas1)
XM3 net4 net4 VSS VSS sg13_hv_nmos w=4.5u l=2u ng=2 m=2
XM4 net1 net1 VSS VSS sg13_hv_nmos w=1u l=3.8u ng=2 m=2
**** begin user architecture code


.param mm_ok=0
.param mc_ok=0
.param temp=27
.param VDD=3.3
.param VSS=0
.control
	save all
	dc temp -40 125 1
	plot i(Vmeas1)
	op
	write op.raw
.endc



.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerRES.lib res_typ


.lib cornerMOShv.lib mos_fs

**** end user architecture code
**.ends
.GLOBAL GND
.end
