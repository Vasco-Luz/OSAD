magic
tech sky130A
magscale 1 2
timestamp 1740493314
<< mvpsubdiff >>
rect -119 1161 -59 1195
rect 1677 1161 1737 1195
rect -119 1135 -85 1161
rect -119 -85 -85 -59
rect 1703 1135 1737 1161
rect 1703 -85 1737 -59
rect -119 -119 -59 -85
rect 1677 -119 1737 -85
<< mvpsubdiffcont >>
rect -59 1161 1677 1195
rect -119 -59 -85 1135
rect 1703 -59 1737 1135
rect -59 -119 1677 -85
<< locali >>
rect -119 1161 -59 1195
rect 1677 1161 1737 1195
rect -119 1135 -85 1161
rect 1703 1135 1737 1161
rect 332 1012 1274 1024
rect 332 978 344 1012
rect 378 978 432 1012
rect 466 978 1274 1012
rect 332 940 1274 978
rect 12 864 98 898
rect 332 864 500 940
rect 12 702 46 864
rect 590 862 758 940
rect 848 864 1016 940
rect 1106 862 1274 940
rect 1514 864 1594 898
rect 1560 776 1594 864
rect -119 -85 -85 -59
rect 12 -85 46 66
rect 270 -85 304 64
rect 786 -85 820 84
rect 1302 -85 1336 68
rect 1560 -85 1594 74
rect 1703 -85 1737 -59
rect -119 -86 -59 -85
rect -120 -119 -59 -86
rect 1677 -119 1737 -85
rect -120 -194 1736 -119
<< viali >>
rect 344 978 378 1012
rect 432 978 466 1012
<< metal1 >>
rect 528 1116 678 1122
rect 528 1062 534 1116
rect 586 1062 620 1116
rect 672 1062 678 1116
rect 528 1056 678 1062
rect 928 1120 1078 1126
rect 928 1066 934 1120
rect 986 1066 1020 1120
rect 1072 1066 1078 1120
rect 928 1060 1078 1066
rect 332 1024 482 1030
rect 332 972 338 1024
rect 390 972 424 1024
rect 476 972 482 1024
rect 332 966 482 972
rect 528 778 562 1056
rect 1044 790 1078 1060
<< via1 >>
rect 534 1062 586 1116
rect 620 1062 672 1116
rect 934 1066 986 1120
rect 1020 1066 1072 1120
rect 338 1012 390 1024
rect 338 978 344 1012
rect 344 978 378 1012
rect 378 978 390 1012
rect 338 972 390 978
rect 424 1012 476 1024
rect 424 978 432 1012
rect 432 978 466 1012
rect 466 978 476 1012
rect 424 972 476 978
<< metal2 >>
rect 528 1116 678 1122
rect 928 1120 1078 1126
rect 928 1116 934 1120
rect 528 1062 534 1116
rect 586 1062 620 1116
rect 672 1066 934 1116
rect 986 1066 1020 1120
rect 1072 1066 1078 1120
rect 672 1062 1078 1066
rect 528 1060 1078 1062
rect 528 1056 678 1060
rect 332 1024 482 1030
rect 132 972 338 1024
rect 390 972 424 1024
rect 476 972 482 1024
rect 332 966 482 972
use sky130_fd_pr__nfet_g5v0d10v5_8F5HCW  sky130_fd_pr__nfet_g5v0d10v5_8F5HCW_0
timestamp 1740484998
transform 1 0 1061 0 1 457
box -287 -457 287 457
use sky130_fd_pr__nfet_g5v0d10v5_8F5HCW  sky130_fd_pr__nfet_g5v0d10v5_8F5HCW_1
timestamp 1740484998
transform 1 0 545 0 1 457
box -287 -457 287 457
use sky130_fd_pr__nfet_g5v0d10v5_JZTFN8  sky130_fd_pr__nfet_g5v0d10v5_JZTFN8_0
timestamp 1740484998
transform 1 0 158 0 1 457
box -158 -457 158 457
use sky130_fd_pr__nfet_g5v0d10v5_JZTFN8  sky130_fd_pr__nfet_g5v0d10v5_JZTFN8_1
timestamp 1740484998
transform 1 0 1448 0 1 457
box -158 -457 158 457
<< labels >>
flabel metal2 152 976 192 1014 0 FreeSans 1600 0 0 0 Ib
port 3 nsew
flabel metal2 796 1074 836 1112 0 FreeSans 1600 0 0 0 VOUT
port 5 nsew
flabel locali 408 -162 482 -136 0 FreeSans 1600 0 0 0 VSS
port 10 nsew
<< end >>
