magic
tech sky130A
magscale 1 2
timestamp 1740409548
<< error_p >>
rect -611 548 611 552
rect -611 -480 -581 548
rect -545 482 545 486
rect -545 -414 -515 482
rect -463 -514 201 -276
rect 515 -414 545 482
rect 581 -480 611 548
rect -209 -530 -53 -514
rect -53 -592 -41 -530
<< nwell >>
rect -581 -514 581 548
rect -209 -592 -53 -530
<< mvpmos >>
rect -487 -414 -287 486
rect -229 -414 -29 486
rect 29 -414 229 486
rect 287 -414 487 486
<< mvpdiff >>
rect -545 474 -487 486
rect -545 -402 -533 474
rect -499 -402 -487 474
rect -545 -414 -487 -402
rect -287 474 -229 486
rect -287 -402 -275 474
rect -241 -402 -229 474
rect -287 -414 -229 -402
rect -29 474 29 486
rect -29 -402 -17 474
rect 17 -402 29 474
rect -29 -414 29 -402
rect 229 474 287 486
rect 229 -402 241 474
rect 275 -402 287 474
rect 229 -414 287 -402
rect 487 474 545 486
rect 487 -402 499 474
rect 533 -402 545 474
rect 487 -414 545 -402
<< mvpdiffc >>
rect -533 -402 -499 474
rect -275 -402 -241 474
rect -17 -402 17 474
rect 241 -402 275 474
rect 499 -402 533 474
<< poly >>
rect -487 486 -287 512
rect -229 486 -29 512
rect 29 486 229 512
rect 287 486 487 512
rect -487 -461 -287 -414
rect -487 -478 -454 -461
rect -470 -495 -454 -478
rect -320 -478 -287 -461
rect -229 -461 -29 -414
rect -229 -478 -196 -461
rect -320 -495 -304 -478
rect -470 -511 -304 -495
rect -212 -495 -196 -478
rect -62 -478 -29 -461
rect 29 -461 229 -414
rect 29 -478 62 -461
rect -62 -495 -46 -478
rect -212 -511 -46 -495
rect 46 -495 62 -478
rect 196 -478 229 -461
rect 287 -461 487 -414
rect 287 -478 320 -461
rect 196 -495 212 -478
rect 46 -511 212 -495
rect 304 -495 320 -478
rect 454 -478 487 -461
rect 454 -495 470 -478
rect 304 -511 470 -495
<< polycont >>
rect -454 -495 -320 -461
rect -196 -495 -62 -461
rect 62 -495 196 -461
rect 320 -495 454 -461
<< locali >>
rect -533 474 -499 622
rect -533 -418 -499 -402
rect -275 474 -241 490
rect -275 -418 -241 -402
rect -17 474 17 666
rect -17 -418 17 -402
rect 241 474 275 490
rect 241 -418 275 -402
rect 499 474 533 628
rect 499 -418 533 -402
rect -471 -461 -45 -460
rect -471 -495 -454 -461
rect -320 -495 -196 -461
rect -62 -495 -45 -461
rect -471 -496 -45 -495
rect 43 -461 471 -460
rect 43 -495 62 -461
rect 196 -495 320 -461
rect 454 -495 471 -461
rect 43 -496 471 -495
<< viali >>
rect -533 -402 -499 474
rect -275 -402 -241 474
rect -17 -402 17 474
rect 241 -402 275 474
rect 499 -402 533 474
rect -454 -495 -320 -461
rect -196 -495 -62 -461
rect 62 -495 196 -461
rect 320 -495 454 -461
<< metal1 >>
rect -277 946 -119 952
rect -277 894 -271 946
rect -219 894 -177 946
rect -125 894 -119 946
rect -277 888 -119 894
rect 119 946 277 952
rect 119 894 125 946
rect 177 894 219 946
rect 271 894 277 946
rect 119 888 277 894
rect -277 486 -241 888
rect 241 486 277 888
rect -539 474 -493 486
rect -539 -402 -533 474
rect -499 -402 -493 474
rect -539 -414 -493 -402
rect -281 474 -235 486
rect -281 -402 -275 474
rect -241 -402 -235 474
rect -281 -414 -235 -402
rect -23 474 23 486
rect -23 -402 -17 474
rect 17 -402 23 474
rect -23 -414 23 -402
rect 235 474 281 486
rect 235 -402 241 474
rect 275 -402 281 474
rect 235 -414 281 -402
rect 493 474 539 486
rect 493 -402 499 474
rect 533 -402 539 474
rect 493 -414 539 -402
rect -466 -461 -308 -455
rect -466 -495 -454 -461
rect -320 -495 -308 -461
rect -466 -501 -308 -495
rect -211 -461 -49 -454
rect -211 -495 -196 -461
rect -62 -495 -49 -461
rect -211 -534 -49 -495
rect 50 -461 208 -455
rect 308 -460 466 -455
rect 50 -495 62 -461
rect 196 -495 208 -461
rect 50 -501 208 -495
rect 293 -461 467 -460
rect 293 -495 320 -461
rect 454 -495 467 -461
rect -211 -586 -203 -534
rect -151 -536 -49 -534
rect -151 -586 -111 -536
rect -211 -588 -111 -586
rect -59 -588 -49 -536
rect -211 -592 -49 -588
rect 293 -538 467 -495
rect 293 -590 299 -538
rect 351 -540 467 -538
rect 351 -590 391 -540
rect 293 -592 391 -590
rect 443 -592 467 -540
rect 293 -596 467 -592
<< via1 >>
rect -271 894 -219 946
rect -177 894 -125 946
rect 125 894 177 946
rect 219 894 271 946
rect -203 -586 -151 -534
rect -111 -588 -59 -536
rect 299 -590 351 -538
rect 391 -592 443 -540
<< metal2 >>
rect -277 946 -119 952
rect 119 946 277 952
rect -277 894 -271 946
rect -219 894 -177 946
rect -125 894 125 946
rect 177 894 219 946
rect 271 894 277 946
rect -277 888 -119 894
rect 119 888 277 894
rect -209 -534 -53 -530
rect -209 -544 -203 -534
rect -645 -572 -203 -544
rect -209 -586 -203 -572
rect -151 -536 -53 -534
rect -151 -586 -111 -536
rect -209 -588 -111 -586
rect -59 -544 -53 -536
rect 293 -538 449 -534
rect 293 -544 299 -538
rect -59 -572 299 -544
rect -59 -588 -53 -572
rect -209 -592 -53 -588
rect 293 -590 299 -572
rect 351 -540 449 -538
rect 351 -590 391 -540
rect 293 -592 391 -590
rect 443 -544 449 -540
rect 443 -572 675 -544
rect 443 -592 449 -572
rect 293 -596 449 -592
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 4.5 l 1 m 1 nf 4 diffcov 100 polycov 80 guard 0 glc 0 grc 0 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 80 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
